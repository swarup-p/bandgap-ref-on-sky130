magic
tech sky130A
timestamp 1615514367
<< nwell >>
rect 0 9600 29104 10000
rect 432 1500 618 9600
<< mvnmos >>
rect 375 1325 675 1425
rect 375 1195 675 1295
<< mvpmos >>
rect 500 1575 550 9575
<< mvndiff >>
rect 340 1416 375 1425
rect 340 1334 349 1416
rect 366 1334 375 1416
rect 340 1325 375 1334
rect 675 1416 710 1425
rect 675 1334 684 1416
rect 701 1334 710 1416
rect 675 1325 710 1334
rect 340 1286 375 1295
rect 340 1204 349 1286
rect 366 1204 375 1286
rect 340 1195 375 1204
rect 675 1286 710 1295
rect 675 1204 684 1286
rect 701 1204 710 1286
rect 675 1195 710 1204
<< mvpdiff >>
rect 465 9300 500 9575
rect 465 9200 474 9300
rect 491 9200 500 9300
rect 465 8800 500 9200
rect 465 8700 474 8800
rect 491 8700 500 8800
rect 465 8300 500 8700
rect 465 8200 474 8300
rect 491 8200 500 8300
rect 465 7800 500 8200
rect 465 7700 474 7800
rect 491 7700 500 7800
rect 465 7300 500 7700
rect 465 7200 474 7300
rect 491 7200 500 7300
rect 465 6800 500 7200
rect 465 6700 474 6800
rect 491 6700 500 6800
rect 465 6300 500 6700
rect 465 6200 474 6300
rect 491 6200 500 6300
rect 465 5800 500 6200
rect 465 5700 474 5800
rect 491 5700 500 5800
rect 465 5300 500 5700
rect 465 5200 474 5300
rect 491 5200 500 5300
rect 465 4800 500 5200
rect 465 4700 474 4800
rect 491 4700 500 4800
rect 465 4300 500 4700
rect 465 4200 474 4300
rect 491 4200 500 4300
rect 465 3800 500 4200
rect 465 3700 474 3800
rect 491 3700 500 3800
rect 465 3300 500 3700
rect 465 3200 474 3300
rect 491 3200 500 3300
rect 465 2800 500 3200
rect 465 2700 474 2800
rect 491 2700 500 2800
rect 465 2300 500 2700
rect 465 2200 474 2300
rect 491 2200 500 2300
rect 465 1800 500 2200
rect 465 1700 474 1800
rect 491 1700 500 1800
rect 465 1575 500 1700
rect 550 9300 585 9575
rect 550 9200 559 9300
rect 576 9200 585 9300
rect 550 8800 585 9200
rect 550 8700 559 8800
rect 576 8700 585 8800
rect 550 8300 585 8700
rect 550 8200 559 8300
rect 576 8200 585 8300
rect 550 7800 585 8200
rect 550 7700 559 7800
rect 576 7700 585 7800
rect 550 7300 585 7700
rect 550 7200 559 7300
rect 576 7200 585 7300
rect 550 6800 585 7200
rect 550 6700 559 6800
rect 576 6700 585 6800
rect 550 6300 585 6700
rect 550 6200 559 6300
rect 576 6200 585 6300
rect 550 5800 585 6200
rect 550 5700 559 5800
rect 576 5700 585 5800
rect 550 5300 585 5700
rect 550 5200 559 5300
rect 576 5200 585 5300
rect 550 4800 585 5200
rect 550 4700 559 4800
rect 576 4700 585 4800
rect 550 4300 585 4700
rect 550 4200 559 4300
rect 576 4200 585 4300
rect 550 3800 585 4200
rect 550 3700 559 3800
rect 576 3700 585 3800
rect 550 3300 585 3700
rect 550 3200 559 3300
rect 576 3200 585 3300
rect 550 2800 585 3200
rect 550 2700 559 2800
rect 576 2700 585 2800
rect 550 2300 585 2700
rect 550 2200 559 2300
rect 576 2200 585 2300
rect 550 1800 585 2200
rect 550 1700 559 1800
rect 576 1700 585 1800
rect 550 1575 585 1700
<< mvndiffc >>
rect 349 1334 366 1416
rect 684 1334 701 1416
rect 349 1204 366 1286
rect 684 1204 701 1286
<< mvpdiffc >>
rect 474 9200 491 9300
rect 474 8700 491 8800
rect 474 8200 491 8300
rect 474 7700 491 7800
rect 474 7200 491 7300
rect 474 6700 491 6800
rect 474 6200 491 6300
rect 474 5700 491 5800
rect 474 5200 491 5300
rect 474 4700 491 4800
rect 474 4200 491 4300
rect 474 3700 491 3800
rect 474 3200 491 3300
rect 474 2700 491 2800
rect 474 2200 491 2300
rect 474 1700 491 1800
rect 559 9200 576 9300
rect 559 8700 576 8800
rect 559 8200 576 8300
rect 559 7700 576 7800
rect 559 7200 576 7300
rect 559 6700 576 6800
rect 559 6200 576 6300
rect 559 5700 576 5800
rect 559 5200 576 5300
rect 559 4700 576 4800
rect 559 4200 576 4300
rect 559 3700 576 3800
rect 559 3200 576 3300
rect 559 2700 576 2800
rect 559 2200 576 2300
rect 559 1700 576 1800
<< mvpsubdiff >>
rect 200 300 28904 390
rect 200 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9920 300
rect 10020 200 10220 300
rect 10320 200 10520 300
rect 10620 200 10820 300
rect 10920 200 11120 300
rect 11220 200 11420 300
rect 11520 200 11720 300
rect 11820 200 12020 300
rect 12120 200 12320 300
rect 12420 200 12620 300
rect 12720 200 12920 300
rect 13020 200 13220 300
rect 13320 200 13520 300
rect 13620 200 13820 300
rect 13920 200 14120 300
rect 14220 200 14420 300
rect 14520 200 14720 300
rect 14820 200 15020 300
rect 15120 200 15320 300
rect 15420 200 15620 300
rect 15720 200 15920 300
rect 16020 200 16220 300
rect 16320 200 16520 300
rect 16620 200 16820 300
rect 16920 200 17120 300
rect 17220 200 17420 300
rect 17520 200 17720 300
rect 17820 200 18020 300
rect 18120 200 18320 300
rect 18420 200 18620 300
rect 18720 200 18920 300
rect 19020 200 19220 300
rect 19320 200 19520 300
rect 19620 200 19820 300
rect 19920 200 20120 300
rect 20220 200 20420 300
rect 20520 200 20720 300
rect 20820 200 21020 300
rect 21120 200 21320 300
rect 21420 200 21620 300
rect 21720 200 21920 300
rect 22020 200 22220 300
rect 22320 200 22520 300
rect 22620 200 22820 300
rect 22920 200 23120 300
rect 23220 200 23420 300
rect 23520 200 23720 300
rect 23820 200 24020 300
rect 24120 200 24320 300
rect 24420 200 24620 300
rect 24720 200 24920 300
rect 25020 200 25220 300
rect 25320 200 25520 300
rect 25620 200 25820 300
rect 25920 200 26120 300
rect 26220 200 26420 300
rect 26520 200 26720 300
rect 26820 200 27020 300
rect 27120 200 27320 300
rect 27420 200 27620 300
rect 27720 200 27920 300
rect 28020 200 28220 300
rect 28320 200 28520 300
rect 28620 200 28904 300
rect 200 110 28904 200
<< mvnsubdiff >>
rect 200 9850 28904 9940
rect 200 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9920 9850
rect 10020 9750 10220 9850
rect 10320 9750 10520 9850
rect 10620 9750 10820 9850
rect 10920 9750 11120 9850
rect 11220 9750 11420 9850
rect 11520 9750 11720 9850
rect 11820 9750 12020 9850
rect 12120 9750 12320 9850
rect 12420 9750 12620 9850
rect 12720 9750 12920 9850
rect 13020 9750 13220 9850
rect 13320 9750 13520 9850
rect 13620 9750 13820 9850
rect 13920 9750 14120 9850
rect 14220 9750 14420 9850
rect 14520 9750 14720 9850
rect 14820 9750 15020 9850
rect 15120 9750 15320 9850
rect 15420 9750 15620 9850
rect 15720 9750 15920 9850
rect 16020 9750 16220 9850
rect 16320 9750 16520 9850
rect 16620 9750 16820 9850
rect 16920 9750 17120 9850
rect 17220 9750 17420 9850
rect 17520 9750 17720 9850
rect 17820 9750 18020 9850
rect 18120 9750 18320 9850
rect 18420 9750 18620 9850
rect 18720 9750 18920 9850
rect 19020 9750 19220 9850
rect 19320 9750 19520 9850
rect 19620 9750 19820 9850
rect 19920 9750 20120 9850
rect 20220 9750 20420 9850
rect 20520 9750 20720 9850
rect 20820 9750 21020 9850
rect 21120 9750 21320 9850
rect 21420 9750 21620 9850
rect 21720 9750 21920 9850
rect 22020 9750 22220 9850
rect 22320 9750 22520 9850
rect 22620 9750 22820 9850
rect 22920 9750 23120 9850
rect 23220 9750 23420 9850
rect 23520 9750 23720 9850
rect 23820 9750 24020 9850
rect 24120 9750 24320 9850
rect 24420 9750 24620 9850
rect 24720 9750 24920 9850
rect 25020 9750 25220 9850
rect 25320 9750 25520 9850
rect 25620 9750 25820 9850
rect 25920 9750 26120 9850
rect 26220 9750 26420 9850
rect 26520 9750 26720 9850
rect 26820 9750 27020 9850
rect 27120 9750 27320 9850
rect 27420 9750 27620 9850
rect 27720 9750 27920 9850
rect 28020 9750 28220 9850
rect 28320 9750 28520 9850
rect 28620 9750 28904 9850
rect 200 9660 28904 9750
<< mvpsubdiffcont >>
rect 320 200 420 300
rect 620 200 720 300
rect 920 200 1020 300
rect 1220 200 1320 300
rect 1520 200 1620 300
rect 1820 200 1920 300
rect 2120 200 2220 300
rect 2420 200 2520 300
rect 2720 200 2820 300
rect 3020 200 3120 300
rect 3320 200 3420 300
rect 3620 200 3720 300
rect 3920 200 4020 300
rect 4220 200 4320 300
rect 4520 200 4620 300
rect 4820 200 4920 300
rect 5120 200 5220 300
rect 5420 200 5520 300
rect 5720 200 5820 300
rect 6020 200 6120 300
rect 6320 200 6420 300
rect 6620 200 6720 300
rect 6920 200 7020 300
rect 7220 200 7320 300
rect 7520 200 7620 300
rect 7820 200 7920 300
rect 8120 200 8220 300
rect 8420 200 8520 300
rect 8720 200 8820 300
rect 9020 200 9120 300
rect 9320 200 9420 300
rect 9620 200 9720 300
rect 9920 200 10020 300
rect 10220 200 10320 300
rect 10520 200 10620 300
rect 10820 200 10920 300
rect 11120 200 11220 300
rect 11420 200 11520 300
rect 11720 200 11820 300
rect 12020 200 12120 300
rect 12320 200 12420 300
rect 12620 200 12720 300
rect 12920 200 13020 300
rect 13220 200 13320 300
rect 13520 200 13620 300
rect 13820 200 13920 300
rect 14120 200 14220 300
rect 14420 200 14520 300
rect 14720 200 14820 300
rect 15020 200 15120 300
rect 15320 200 15420 300
rect 15620 200 15720 300
rect 15920 200 16020 300
rect 16220 200 16320 300
rect 16520 200 16620 300
rect 16820 200 16920 300
rect 17120 200 17220 300
rect 17420 200 17520 300
rect 17720 200 17820 300
rect 18020 200 18120 300
rect 18320 200 18420 300
rect 18620 200 18720 300
rect 18920 200 19020 300
rect 19220 200 19320 300
rect 19520 200 19620 300
rect 19820 200 19920 300
rect 20120 200 20220 300
rect 20420 200 20520 300
rect 20720 200 20820 300
rect 21020 200 21120 300
rect 21320 200 21420 300
rect 21620 200 21720 300
rect 21920 200 22020 300
rect 22220 200 22320 300
rect 22520 200 22620 300
rect 22820 200 22920 300
rect 23120 200 23220 300
rect 23420 200 23520 300
rect 23720 200 23820 300
rect 24020 200 24120 300
rect 24320 200 24420 300
rect 24620 200 24720 300
rect 24920 200 25020 300
rect 25220 200 25320 300
rect 25520 200 25620 300
rect 25820 200 25920 300
rect 26120 200 26220 300
rect 26420 200 26520 300
rect 26720 200 26820 300
rect 27020 200 27120 300
rect 27320 200 27420 300
rect 27620 200 27720 300
rect 27920 200 28020 300
rect 28220 200 28320 300
rect 28520 200 28620 300
<< mvnsubdiffcont >>
rect 320 9750 420 9850
rect 620 9750 720 9850
rect 920 9750 1020 9850
rect 1220 9750 1320 9850
rect 1520 9750 1620 9850
rect 1820 9750 1920 9850
rect 2120 9750 2220 9850
rect 2420 9750 2520 9850
rect 2720 9750 2820 9850
rect 3020 9750 3120 9850
rect 3320 9750 3420 9850
rect 3620 9750 3720 9850
rect 3920 9750 4020 9850
rect 4220 9750 4320 9850
rect 4520 9750 4620 9850
rect 4820 9750 4920 9850
rect 5120 9750 5220 9850
rect 5420 9750 5520 9850
rect 5720 9750 5820 9850
rect 6020 9750 6120 9850
rect 6320 9750 6420 9850
rect 6620 9750 6720 9850
rect 6920 9750 7020 9850
rect 7220 9750 7320 9850
rect 7520 9750 7620 9850
rect 7820 9750 7920 9850
rect 8120 9750 8220 9850
rect 8420 9750 8520 9850
rect 8720 9750 8820 9850
rect 9020 9750 9120 9850
rect 9320 9750 9420 9850
rect 9620 9750 9720 9850
rect 9920 9750 10020 9850
rect 10220 9750 10320 9850
rect 10520 9750 10620 9850
rect 10820 9750 10920 9850
rect 11120 9750 11220 9850
rect 11420 9750 11520 9850
rect 11720 9750 11820 9850
rect 12020 9750 12120 9850
rect 12320 9750 12420 9850
rect 12620 9750 12720 9850
rect 12920 9750 13020 9850
rect 13220 9750 13320 9850
rect 13520 9750 13620 9850
rect 13820 9750 13920 9850
rect 14120 9750 14220 9850
rect 14420 9750 14520 9850
rect 14720 9750 14820 9850
rect 15020 9750 15120 9850
rect 15320 9750 15420 9850
rect 15620 9750 15720 9850
rect 15920 9750 16020 9850
rect 16220 9750 16320 9850
rect 16520 9750 16620 9850
rect 16820 9750 16920 9850
rect 17120 9750 17220 9850
rect 17420 9750 17520 9850
rect 17720 9750 17820 9850
rect 18020 9750 18120 9850
rect 18320 9750 18420 9850
rect 18620 9750 18720 9850
rect 18920 9750 19020 9850
rect 19220 9750 19320 9850
rect 19520 9750 19620 9850
rect 19820 9750 19920 9850
rect 20120 9750 20220 9850
rect 20420 9750 20520 9850
rect 20720 9750 20820 9850
rect 21020 9750 21120 9850
rect 21320 9750 21420 9850
rect 21620 9750 21720 9850
rect 21920 9750 22020 9850
rect 22220 9750 22320 9850
rect 22520 9750 22620 9850
rect 22820 9750 22920 9850
rect 23120 9750 23220 9850
rect 23420 9750 23520 9850
rect 23720 9750 23820 9850
rect 24020 9750 24120 9850
rect 24320 9750 24420 9850
rect 24620 9750 24720 9850
rect 24920 9750 25020 9850
rect 25220 9750 25320 9850
rect 25520 9750 25620 9850
rect 25820 9750 25920 9850
rect 26120 9750 26220 9850
rect 26420 9750 26520 9850
rect 26720 9750 26820 9850
rect 27020 9750 27120 9850
rect 27320 9750 27420 9850
rect 27620 9750 27720 9850
rect 27920 9750 28020 9850
rect 28220 9750 28320 9850
rect 28520 9750 28620 9850
<< poly >>
rect 500 9575 550 9600
rect 500 1542 550 1575
rect 500 1510 516 1542
rect 534 1510 550 1542
rect 500 1500 550 1510
rect 375 1478 675 1500
rect 375 1446 516 1478
rect 534 1446 675 1478
rect 375 1425 675 1446
rect 375 1295 675 1325
rect 375 1175 675 1195
rect 375 1143 516 1175
rect 534 1143 675 1175
rect 375 1135 675 1143
<< polycont >>
rect 516 1510 534 1542
rect 516 1446 534 1478
rect 516 1143 534 1175
<< locali >>
rect 100 9850 29004 9940
rect 100 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9920 9850
rect 10020 9750 10220 9850
rect 10320 9750 10520 9850
rect 10620 9750 10820 9850
rect 10920 9750 11120 9850
rect 11220 9750 11420 9850
rect 11520 9750 11720 9850
rect 11820 9750 12020 9850
rect 12120 9750 12320 9850
rect 12420 9750 12620 9850
rect 12720 9750 12920 9850
rect 13020 9750 13220 9850
rect 13320 9750 13520 9850
rect 13620 9750 13820 9850
rect 13920 9750 14120 9850
rect 14220 9750 14420 9850
rect 14520 9750 14720 9850
rect 14820 9750 15020 9850
rect 15120 9750 15320 9850
rect 15420 9750 15620 9850
rect 15720 9750 15920 9850
rect 16020 9750 16220 9850
rect 16320 9750 16520 9850
rect 16620 9750 16820 9850
rect 16920 9750 17120 9850
rect 17220 9750 17420 9850
rect 17520 9750 17720 9850
rect 17820 9750 18020 9850
rect 18120 9750 18320 9850
rect 18420 9750 18620 9850
rect 18720 9750 18920 9850
rect 19020 9750 19220 9850
rect 19320 9750 19520 9850
rect 19620 9750 19820 9850
rect 19920 9750 20120 9850
rect 20220 9750 20420 9850
rect 20520 9750 20720 9850
rect 20820 9750 21020 9850
rect 21120 9750 21320 9850
rect 21420 9750 21620 9850
rect 21720 9750 21920 9850
rect 22020 9750 22220 9850
rect 22320 9750 22520 9850
rect 22620 9750 22820 9850
rect 22920 9750 23120 9850
rect 23220 9750 23420 9850
rect 23520 9750 23720 9850
rect 23820 9750 24020 9850
rect 24120 9750 24320 9850
rect 24420 9750 24620 9850
rect 24720 9750 24920 9850
rect 25020 9750 25220 9850
rect 25320 9750 25520 9850
rect 25620 9750 25820 9850
rect 25920 9750 26120 9850
rect 26220 9750 26420 9850
rect 26520 9750 26720 9850
rect 26820 9750 27020 9850
rect 27120 9750 27320 9850
rect 27420 9750 27620 9850
rect 27720 9750 27920 9850
rect 28020 9750 28220 9850
rect 28320 9750 28520 9850
rect 28620 9750 29004 9850
rect 100 9660 29004 9750
rect 474 9300 491 9660
rect 474 8800 491 9200
rect 474 8300 491 8700
rect 474 7800 491 8200
rect 474 7300 491 7700
rect 474 6800 491 7200
rect 474 6300 491 6700
rect 474 5800 491 6200
rect 474 5300 491 5700
rect 474 4800 491 5200
rect 474 4300 491 4700
rect 474 3800 491 4200
rect 474 3300 491 3700
rect 474 2800 491 3200
rect 474 2300 491 2700
rect 474 1800 491 2200
rect 474 1575 491 1700
rect 559 9300 576 9575
rect 559 8800 576 9200
rect 559 8300 576 8700
rect 559 7800 576 8200
rect 559 7300 576 7700
rect 559 6800 576 7200
rect 559 6300 576 6700
rect 559 5800 576 6200
rect 559 5300 576 5700
rect 559 4800 576 5200
rect 559 4300 576 4700
rect 559 3800 576 4200
rect 559 3300 576 3700
rect 559 2800 576 3200
rect 559 2300 576 2700
rect 559 1800 576 2200
rect 559 1545 576 1700
rect 506 1542 576 1545
rect 506 1510 516 1542
rect 534 1510 576 1542
rect 506 1508 576 1510
rect 559 1480 576 1508
rect 506 1478 576 1480
rect 506 1446 516 1478
rect 534 1446 576 1478
rect 506 1444 576 1446
rect 349 1416 366 1425
rect 349 1286 366 1334
rect 349 390 366 1204
rect 684 1416 701 1425
rect 684 1286 701 1334
rect 684 1178 701 1204
rect 506 1175 701 1178
rect 506 1143 516 1175
rect 534 1143 701 1175
rect 506 1141 701 1143
rect 100 300 29004 390
rect 100 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9920 300
rect 10020 200 10220 300
rect 10320 200 10520 300
rect 10620 200 10820 300
rect 10920 200 11120 300
rect 11220 200 11420 300
rect 11520 200 11720 300
rect 11820 200 12020 300
rect 12120 200 12320 300
rect 12420 200 12620 300
rect 12720 200 12920 300
rect 13020 200 13220 300
rect 13320 200 13520 300
rect 13620 200 13820 300
rect 13920 200 14120 300
rect 14220 200 14420 300
rect 14520 200 14720 300
rect 14820 200 15020 300
rect 15120 200 15320 300
rect 15420 200 15620 300
rect 15720 200 15920 300
rect 16020 200 16220 300
rect 16320 200 16520 300
rect 16620 200 16820 300
rect 16920 200 17120 300
rect 17220 200 17420 300
rect 17520 200 17720 300
rect 17820 200 18020 300
rect 18120 200 18320 300
rect 18420 200 18620 300
rect 18720 200 18920 300
rect 19020 200 19220 300
rect 19320 200 19520 300
rect 19620 200 19820 300
rect 19920 200 20120 300
rect 20220 200 20420 300
rect 20520 200 20720 300
rect 20820 200 21020 300
rect 21120 200 21320 300
rect 21420 200 21620 300
rect 21720 200 21920 300
rect 22020 200 22220 300
rect 22320 200 22520 300
rect 22620 200 22820 300
rect 22920 200 23120 300
rect 23220 200 23420 300
rect 23520 200 23720 300
rect 23820 200 24020 300
rect 24120 200 24320 300
rect 24420 200 24620 300
rect 24720 200 24920 300
rect 25020 200 25220 300
rect 25320 200 25520 300
rect 25620 200 25820 300
rect 25920 200 26120 300
rect 26220 200 26420 300
rect 26520 200 26720 300
rect 26820 200 27020 300
rect 27120 200 27320 300
rect 27420 200 27620 300
rect 27720 200 27920 300
rect 28020 200 28220 300
rect 28320 200 28520 300
rect 28620 200 29004 300
rect 100 110 29004 200
<< metal1 >>
rect 0 9650 29104 9950
rect 0 0 29104 500
<< end >>
