magic
tech sky130A
magscale 1 2
timestamp 1616542016
<< nwell >>
rect -706 19202 9000 20000
rect -706 17320 -396 19202
rect 0 19200 9000 19202
rect 1536 15050 5860 19200
<< mvpsubdiff >>
rect 400 2380 8600 2560
rect 400 2180 640 2380
rect 840 2180 1240 2380
rect 1440 2180 1840 2380
rect 2040 2180 2440 2380
rect 2640 2180 3040 2380
rect 3240 2180 3640 2380
rect 3840 2180 4240 2380
rect 4440 2180 4840 2380
rect 5040 2180 5440 2380
rect 5640 2180 6040 2380
rect 6240 2180 6640 2380
rect 6840 2180 7240 2380
rect 7440 2180 7840 2380
rect 8040 2180 8600 2380
rect 400 2000 8600 2180
<< mvnsubdiff >>
rect 400 19700 8600 19880
rect 400 19500 640 19700
rect 840 19500 1240 19700
rect 1440 19500 1840 19700
rect 2040 19500 2440 19700
rect 2640 19500 3040 19700
rect 3240 19500 3640 19700
rect 3840 19500 4240 19700
rect 4440 19500 4840 19700
rect 5040 19500 5440 19700
rect 5640 19500 6040 19700
rect 6240 19500 6640 19700
rect 6840 19500 7240 19700
rect 7440 19500 7840 19700
rect 8040 19500 8600 19700
rect 400 19320 8600 19500
<< mvpsubdiffcont >>
rect 640 2180 840 2380
rect 1240 2180 1440 2380
rect 1840 2180 2040 2380
rect 2440 2180 2640 2380
rect 3040 2180 3240 2380
rect 3640 2180 3840 2380
rect 4240 2180 4440 2380
rect 4840 2180 5040 2380
rect 5440 2180 5640 2380
rect 6040 2180 6240 2380
rect 6640 2180 6840 2380
rect 7240 2180 7440 2380
rect 7840 2180 8040 2380
<< mvnsubdiffcont >>
rect 640 19500 840 19700
rect 1240 19500 1440 19700
rect 1840 19500 2040 19700
rect 2440 19500 2640 19700
rect 3040 19500 3240 19700
rect 3640 19500 3840 19700
rect 4240 19500 4440 19700
rect 4840 19500 5040 19700
rect 5440 19500 5640 19700
rect 6040 19500 6240 19700
rect 6640 19500 6840 19700
rect 7240 19500 7440 19700
rect 7840 19500 8040 19700
<< poly >>
rect 2672 18230 3198 19170
rect 2672 18180 3146 18230
rect 3180 18180 3198 18230
rect 2672 18170 3198 18180
rect 4198 18170 4724 19170
rect 2672 13840 3198 14840
rect 2672 9540 3198 10540
rect 4198 9540 4724 10540
<< polycont >>
rect 1688 18204 1738 18238
rect 3146 18180 3180 18230
rect 1040 15068 1108 15102
rect 356 14272 556 14306
rect 1692 14272 1742 14306
rect 1692 13954 1742 13988
rect -450 5288 -416 5356
<< xpolycontact >>
rect 6360 15574 6430 16006
rect 6042 9222 6112 9654
rect 6042 7040 6112 7472
rect 6360 7040 6430 7472
rect 6678 15574 6748 16006
rect 6678 7040 6748 7472
<< xpolyres >>
rect 6042 7472 6112 9222
rect 6360 7472 6430 15574
rect 6678 7472 6748 15574
<< locali >>
rect 200 19700 8800 19880
rect 200 19582 640 19700
rect -566 19548 640 19582
rect -566 17308 -532 19548
rect 200 19500 640 19548
rect 840 19500 1240 19700
rect 1440 19500 1840 19700
rect 2040 19500 2440 19700
rect 2640 19500 3040 19700
rect 3240 19500 3640 19700
rect 3840 19500 4240 19700
rect 4440 19500 4840 19700
rect 5040 19500 5440 19700
rect 5640 19500 6040 19700
rect 6240 19500 6640 19700
rect 6840 19500 7240 19700
rect 7440 19500 7840 19700
rect 8040 19500 8800 19700
rect 200 19320 8800 19500
rect 918 18204 1688 18238
rect 1738 18204 1754 18238
rect 918 15752 952 18204
rect 2690 18120 2724 19320
rect 3146 18230 3180 18246
rect 3146 18120 3180 18180
rect 4216 18120 4250 19320
rect 5742 18120 5776 19320
rect 6358 16006 6432 16008
rect 6358 15574 6360 16006
rect 6430 15804 6432 16006
rect 6676 16006 6750 16008
rect 6676 15804 6678 16006
rect 6430 15770 6678 15804
rect 6430 15574 6432 15770
rect 6358 15572 6432 15574
rect 6676 15574 6678 15770
rect 6748 15574 6750 16006
rect 6676 15572 6750 15574
rect -308 15068 1040 15102
rect 1108 15068 1124 15102
rect -450 5356 -416 5372
rect -450 5238 -416 5288
rect -308 5238 -274 15068
rect 1188 14578 1222 15152
rect 1620 15096 1654 15120
rect 1620 15040 1654 15046
rect 3146 15096 3180 15120
rect 3146 15040 3180 15046
rect 4672 15096 4706 15120
rect 4672 15040 4706 15046
rect 1188 14512 1222 14528
rect 340 14272 356 14306
rect 556 14272 1692 14306
rect 1742 14272 1768 14306
rect 1620 13954 1692 13988
rect 1742 13954 1758 13988
rect 1188 13912 1222 13918
rect -502 5204 -148 5238
rect 1088 5176 1122 5222
rect 1188 5176 1222 13862
rect 1620 13862 1654 13954
rect 1620 13790 1654 13812
rect 3146 13862 3180 13950
rect 3146 13790 3180 13812
rect 2690 10766 2724 10790
rect 2690 10710 2724 10716
rect 4216 10766 4250 10790
rect 4216 10710 4250 10716
rect 3146 9656 6114 9690
rect 2690 9564 2724 9570
rect 2690 9490 2724 9514
rect 3146 9490 3180 9656
rect 6040 9654 6114 9656
rect 4216 9564 4250 9570
rect 4216 9490 4250 9514
rect 4672 9564 4706 9570
rect 4672 9490 4706 9514
rect 6040 9222 6042 9654
rect 6112 9222 6114 9654
rect 6040 9220 6114 9222
rect 6040 7472 6114 7474
rect 1620 7066 1654 7090
rect 1620 7010 1654 7016
rect 5742 7022 5776 7090
rect 5742 6960 5776 6972
rect 6040 7040 6042 7472
rect 6112 7040 6114 7472
rect 6040 6932 6114 7040
rect 6358 7472 6432 7474
rect 6358 7040 6360 7472
rect 6430 7040 6432 7472
rect 6358 7022 6432 7040
rect 6358 6972 6378 7022
rect 6412 6972 6432 7022
rect 6358 6960 6432 6972
rect 6676 7472 6750 7474
rect 6676 7040 6678 7472
rect 6748 7040 6750 7472
rect 6676 7020 6750 7040
rect 6676 6970 6696 7020
rect 6730 6970 6750 7020
rect 6676 6960 6750 6970
rect 6040 6882 6060 6932
rect 6094 6882 6114 6932
rect 6040 6872 6114 6882
rect 1600 6036 1672 6100
rect 2398 6036 2470 6100
rect 3196 6036 3268 6100
rect 3994 6036 4066 6100
rect 4792 6036 4864 6100
rect 1264 5916 5200 5936
rect 1264 5882 5354 5916
rect 1264 5864 5200 5882
rect 1600 5220 1672 5284
rect 2398 5220 2470 5284
rect 3196 5220 3268 5284
rect 3994 5220 4066 5284
rect 4792 5220 4864 5284
rect 1088 5142 1222 5176
rect 1188 2560 1222 5142
rect 5320 2560 5354 5882
rect 200 2380 8800 2560
rect 200 2180 640 2380
rect 840 2180 1240 2380
rect 1440 2180 1840 2380
rect 2040 2180 2440 2380
rect 2640 2180 3040 2380
rect 3240 2180 3640 2380
rect 3840 2180 4240 2380
rect 4440 2180 4840 2380
rect 5040 2180 5440 2380
rect 5640 2180 6040 2380
rect 6240 2180 6640 2380
rect 6840 2180 7240 2380
rect 7440 2180 7840 2380
rect 8040 2180 8800 2380
rect 200 2000 8800 2180
<< viali >>
rect 640 19500 840 19700
rect 1240 19500 1440 19700
rect 1840 19500 2040 19700
rect 2440 19500 2640 19700
rect 3040 19500 3240 19700
rect 3640 19500 3840 19700
rect 4240 19500 4440 19700
rect 4840 19500 5040 19700
rect 5440 19500 5640 19700
rect 6040 19500 6240 19700
rect 6640 19500 6840 19700
rect 7240 19500 7440 19700
rect 7840 19500 8040 19700
rect 1620 15046 1654 15096
rect 3146 15046 3180 15096
rect 4672 15046 4706 15096
rect 1188 14528 1222 14578
rect 1188 13862 1222 13912
rect 1620 13812 1654 13862
rect 3146 13812 3180 13862
rect 2690 10716 2724 10766
rect 4216 10716 4250 10766
rect 2690 9514 2724 9564
rect 4216 9514 4250 9564
rect 4672 9514 4706 9564
rect 1620 7016 1654 7066
rect 5742 6972 5776 7022
rect 6378 6972 6412 7022
rect 6696 6970 6730 7020
rect 6060 6882 6094 6932
rect 640 2180 840 2380
rect 1240 2180 1440 2380
rect 1840 2180 2040 2380
rect 2440 2180 2640 2380
rect 3040 2180 3240 2380
rect 3640 2180 3840 2380
rect 4240 2180 4440 2380
rect 4840 2180 5040 2380
rect 5440 2180 5640 2380
rect 6040 2180 6240 2380
rect 6640 2180 6840 2380
rect 7240 2180 7440 2380
rect 7840 2180 8040 2380
<< metal1 >>
rect 0 19700 9000 19900
rect 0 19500 640 19700
rect 840 19500 1240 19700
rect 1440 19500 1840 19700
rect 2040 19500 2440 19700
rect 2640 19500 3040 19700
rect 3240 19500 3640 19700
rect 3840 19500 4240 19700
rect 4440 19500 4840 19700
rect 5040 19500 5440 19700
rect 5640 19500 6040 19700
rect 6240 19500 6640 19700
rect 6840 19500 7240 19700
rect 7440 19500 7840 19700
rect 8040 19500 9000 19700
rect 0 19300 9000 19500
rect 1606 15096 1666 15110
rect 1606 15046 1620 15096
rect 1654 15046 1666 15096
rect 1174 14578 1234 14590
rect 1174 14528 1188 14578
rect 1222 14528 1234 14578
rect 1174 13912 1234 14528
rect 1174 13862 1188 13912
rect 1222 13862 1234 13912
rect 1174 13848 1234 13862
rect 1606 13862 1666 15046
rect 1606 13812 1620 13862
rect 1654 13812 1666 13862
rect 1606 13800 1666 13812
rect 3132 15096 3192 15110
rect 3132 15046 3146 15096
rect 3180 15046 3192 15096
rect 3132 13862 3192 15046
rect 3132 13812 3146 13862
rect 3180 13812 3192 13862
rect 3132 13800 3192 13812
rect 4658 15096 4718 15110
rect 4658 15046 4672 15096
rect 4706 15046 4718 15096
rect 2678 10766 2738 10780
rect 2678 10716 2690 10766
rect 2724 10716 2738 10766
rect 2678 9564 2738 10716
rect 2678 9514 2690 9564
rect 2724 9514 2738 9564
rect 2678 9500 2738 9514
rect 4204 10766 4264 10780
rect 4204 10716 4216 10766
rect 4250 10716 4264 10766
rect 4204 9564 4264 10716
rect 4204 9514 4216 9564
rect 4250 9514 4264 9564
rect 4204 9500 4264 9514
rect 4658 9564 4718 15046
rect 4658 9514 4672 9564
rect 4706 9514 4718 9564
rect 4658 9500 4718 9514
rect 1606 7066 1666 7080
rect 1606 7016 1620 7066
rect 1654 7016 1666 7066
rect 1606 6390 1666 7016
rect 5730 7022 6424 7028
rect 5730 6972 5742 7022
rect 5776 6972 6378 7022
rect 6412 6972 6424 7022
rect 5730 6966 6424 6972
rect 6682 7020 6742 7032
rect 6682 6970 6696 7020
rect 6730 6970 6742 7020
rect 3094 6932 6114 6938
rect 3094 6882 6060 6932
rect 6094 6882 6114 6932
rect 3094 6876 6114 6882
rect 3094 6790 3154 6876
rect 1978 6730 4858 6790
rect 1978 5522 2038 6730
rect 2404 6390 2464 6730
rect 2776 5522 2836 6730
rect 3202 6390 3262 6730
rect 3574 5522 3634 6730
rect 4000 6390 4060 6730
rect 4372 5522 4432 6730
rect 4798 6390 4858 6730
rect 6682 5522 6742 6970
rect 1718 5462 2038 5522
rect 2516 5462 2836 5522
rect 3314 5462 3634 5522
rect 4112 5462 4432 5522
rect 4910 5462 6742 5522
rect 0 2380 9000 2780
rect 0 2180 640 2380
rect 840 2180 1240 2380
rect 1440 2180 1840 2380
rect 2040 2180 2440 2380
rect 2640 2180 3040 2380
rect 3240 2180 3640 2380
rect 3840 2180 4240 2380
rect 4440 2180 4840 2380
rect 5040 2180 5440 2380
rect 5640 2180 6040 2380
rect 6240 2180 6640 2380
rect 6840 2180 7240 2380
rect 7440 2180 7840 2380
rect 8040 2180 9000 2380
rect 0 1780 9000 2180
use sc_nmos  sc_nmos_2
timestamp 1616174596
transform 1 0 520 0 1 13950
box 380 1100 720 1904
use sc_nmos_change  sc_nmos_change_0
timestamp 1616538694
transform 1 0 -580 0 1 4020
box 380 1100 1720 10304
use cm_nmos  cm_nmos_1
timestamp 1616067151
transform 1 0 1672 0 1 10740
box -70 0 1070 4100
use en_nmos  en_nmos_0
timestamp 1616065709
transform 1 0 1672 0 1 7040
box -70 0 1070 3500
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 1238 0 1 5094
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 1238 0 1 5910
box 26 26 770 795
use cm_pmos  cm_pmos_0
timestamp 1616078161
transform 1 0 1672 0 1 15070
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 2036 0 1 5094
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 2036 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 2834 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 2834 0 1 5094
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 3632 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 3632 0 1 5094
box 26 26 770 795
use en_nmos  en_nmos_1
timestamp 1616065709
transform 1 0 3198 0 1 7040
box -70 0 1070 3500
use cm_nmos  cm_nmos_0
timestamp 1616067151
transform 1 0 3198 0 1 10740
box -70 0 1070 4100
use cm_pmos  cm_pmos_1
timestamp 1616078161
transform 1 0 3198 0 1 15070
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 4430 0 1 5094
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 4430 0 1 5910
box 26 26 770 795
use en_nmos  en_nmos_2
timestamp 1616065709
transform 1 0 4724 0 1 7040
box -70 0 1070 3500
use cm_pmos  cm_pmos_2
timestamp 1616078161
transform 1 0 4724 0 1 15070
box -136 -20 1136 4100
use sc_pmos  sc_pmos_0
timestamp 1616540248
transform 1 0 -1100 0 1 2192
box 400 2928 700 15200
<< labels >>
flabel locali s 218 19646 640 19934 0 FreeSans 1600 0 0 0 VDD
flabel locali s 238 2338 628 2548 0 FreeSans 1600 0 0 0 GND
flabel poly s 2754 10146 3176 10506 0 FreeSans 1600 0 0 0 en
flabel locali s 6422 6962 6432 6966 0 FreeSans 400 0 0 0 Vbgp
flabel metal1 s 5896 6886 5954 6902 0 FreeSans 400 0 0 0 A
flabel locali s 5900 9662 5958 9678 0 FreeSans 400 0 0 0 B
flabel metal1 s 4216 10642 4274 10658 0 FreeSans 400 0 0 0 C
flabel metal1 s 3168 14956 3226 14972 0 FreeSans 400 0 0 0 D
flabel metal1 s 4694 14940 4708 14960 0 FreeSans 400 0 0 0 E
flabel metal1 s 1646 6976 1660 6996 0 FreeSans 400 0 0 0 F
flabel metal1 s 2704 10660 2718 10680 0 FreeSans 400 0 0 0 G
flabel locali s 6534 15786 6548 15806 0 FreeSans 400 0 0 0 H
flabel metal1 s 6702 6792 6716 6812 0 FreeSans 400 0 0 0 J
flabel locali s 1126 18222 1146 18232 0 FreeSans 1600 0 0 0 VbiasP
flabel locali s 1482 14286 1500 14294 0 FreeSans 800 0 0 0 VbiasN
flabel locali s -378 5220 -360 5228 0 FreeSans 800 0 0 0 I
<< end >>
