magic
tech sky130A
timestamp 1616000842
<< xpolycontact >>
rect 0 489 216 524
rect 8318 489 8534 524
rect 0 326 216 361
rect 492 326 708 361
rect 0 163 216 198
rect 285 163 501 198
rect 0 0 216 35
rect 251 0 467 35
<< xpolyres >>
rect 216 489 8318 524
rect 216 326 492 361
rect 216 163 285 198
rect 216 0 251 35
<< locali >>
rect 0 524 216 528
rect 0 485 216 489
rect 8318 524 8534 528
rect 8318 485 8534 489
rect 0 361 216 363
rect 0 322 216 326
rect 492 361 708 365
rect 492 322 708 326
rect 100 202 117 322
rect 0 198 216 202
rect 0 159 216 163
rect 285 198 501 202
rect 285 159 501 163
rect 0 35 216 39
rect 0 -4 216 0
rect 251 35 467 39
rect 251 -4 467 0
<< end >>
