* SPICE3 file created from bgr_a2.ext - technology: sky130A

.option scale=10000u

X0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/a_330_330# sky130_fd_pr__pnp_05v5_W3p40L3p40_0/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# sky130_fd_pr__pnp_05v0 area=8
X1 m1_2049_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_1/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# sky130_fd_pr__pnp_05v0 area=524287
X2 m1_2793_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_2/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# sky130_fd_pr__pnp_05v0 area=-5.44224e+08
X3 m1_3537_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_3/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# sky130_fd_pr__pnp_05v0 area=97
X4 m1_4281_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_4/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X5 m1_4183_2199# sky130_fd_pr__pnp_05v5_W3p40L3p40_5/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# sky130_fd_pr__pnp_05v0 area=8
X6 m1_3439_2199# sky130_fd_pr__pnp_05v5_W3p40L3p40_6/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X7 m1_2695_2199# sky130_fd_pr__pnp_05v5_W3p40L3p40_7/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# sky130_fd_pr__pnp_05v0 area=8
X8 m1_1951_2199# sky130_fd_pr__pnp_05v5_W3p40L3p40_8/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X9 a_225_550# a_325_1028# w_0_9600# w_0_9600# sky130_fd_pr__pfet_g5v0d10v5 w=1500 l=500
X10 a_325_1028# a_190_601# a_190_1028# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=300 l=100
X11 a_325_1028# a_325_1028# w_0_9600# w_0_9600# sky130_fd_pr__pfet_g5v0d10v5 w=1500 l=500
X12 a_2840_4177# a_325_1028# w_0_9600# w_0_9600# sky130_fd_pr__pfet_g5v0d10v5 w=1500 l=500
X13 a_225_550# a_225_550# a_733_4177# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=1500 l=500
X14 a_250_9532# a_190_601# a_190_601# w_0_9600# sky130_fd_pr__pfet_g5v0d10v5 w=50 l=8000
X15 a_325_1028# a_225_550# a_1519_4177# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=1500 l=500
X16 a_190_1028# a_225_550# a_190_601# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=300 l=100
X17 a_1268_4177# a_768_4126# a_733_4177# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=1200 l=500
X18 a_2054_4177# a_1554_4126# a_1519_4177# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=1200 l=500
X19 a_2840_4177# a_2340_4126# a_2305_4177# a_200_110# sky130_fd_pr__nfet_g5v0d10v5 w=1200 l=500
C0 a_190_601# a_225_550# 2.14fF
C1 m1_2793_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_2/w_153_153# 0.55fF
C2 a_190_601# a_325_1028# 4.29fF
C3 a_733_4177# a_225_550# 0.00fF
C4 a_1554_4126# a_1519_4177# 0.03fF
C5 m1_4183_2199# sky130_fd_pr__pnp_05v5_W3p40L3p40_5/w_153_153# 0.32fF
C6 a_250_9532# w_0_9600# 0.02fF
C7 a_768_4126# a_733_4177# 0.03fF
C8 sky130_fd_pr__pnp_05v5_W3p40L3p40_6/w_153_153# m1_3439_2199# 0.55fF
C9 a_325_1028# a_225_550# 7.11fF
C10 sky130_fd_pr__pnp_05v5_W3p40L3p40_7/w_153_153# m1_2695_2199# 0.55fF
C11 sky130_fd_pr__pnp_05v5_W3p40L3p40_8/w_153_153# m1_1951_2199# 0.55fF
C12 w_0_9600# a_2840_4177# 0.00fF
C13 a_190_601# w_0_9600# 0.01fF
C14 m1_2049_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_1/w_153_153# 0.55fF
C15 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/w_153_153# sky130_fd_pr__pnp_05v5_W3p40L3p40_0/a_330_330# 0.36fF
C16 m1_4281_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_4/w_153_153# 0.55fF
C17 a_190_601# a_190_1028# 0.61fF
C18 w_0_9600# a_225_550# 0.01fF
C19 w_0_9600# m1_0_9650# 39.04fF
C20 a_325_1028# w_0_9600# 0.07fF
C21 a_1519_4177# a_225_550# 0.03fF
C22 a_225_550# a_190_1028# 0.24fF
C23 m1_3537_1357# sky130_fd_pr__pnp_05v5_W3p40L3p40_3/w_153_153# 0.55fF
C24 a_325_1028# a_190_1028# 0.12fF
C25 m1_0_9650# a_200_110# 8.43fF **FLOATING
C26 a_190_1028# a_200_110# 53.43fF
C27 a_2305_4177# a_200_110# 0.02fF
C28 a_2054_4177# a_200_110# 0.02fF
C29 a_1268_4177# a_200_110# 0.02fF
C30 a_2340_4126# a_200_110# 1.22fF
C31 a_1554_4126# a_200_110# 1.21fF
C32 a_768_4126# a_200_110# 1.21fF
C33 a_1519_4177# a_200_110# 0.49fF
C34 a_733_4177# a_200_110# 0.49fF
C35 a_2840_4177# a_200_110# 3.72fF
C36 a_225_550# a_200_110# 14.70fF
C37 a_325_1028# a_200_110# 15.24fF
C38 a_190_601# a_200_110# 18.97fF
C39 a_250_9532# a_200_110# 0.02fF
C40 w_0_9600# a_200_110# 120.19fF
C41 m1_1951_2199# a_200_110# 0.30fF
C42 sky130_fd_pr__pnp_05v5_W3p40L3p40_8/w_153_153# a_200_110# 2.41fF
C43 m1_2695_2199# a_200_110# 0.30fF
C44 sky130_fd_pr__pnp_05v5_W3p40L3p40_7/w_153_153# a_200_110# 2.41fF
C45 m1_3439_2199# a_200_110# 0.80fF
C46 sky130_fd_pr__pnp_05v5_W3p40L3p40_6/w_153_153# a_200_110# 2.41fF
C47 m1_4183_2199# a_200_110# 0.54fF
C48 sky130_fd_pr__pnp_05v5_W3p40L3p40_5/w_153_153# a_200_110# 2.41fF
C49 sky130_fd_pr__pnp_05v5_W3p40L3p40_4/w_153_153# a_200_110# 2.41fF
C50 m1_3537_1357# a_200_110# 0.00fF
C51 sky130_fd_pr__pnp_05v5_W3p40L3p40_3/w_153_153# a_200_110# 2.41fF
C52 sky130_fd_pr__pnp_05v5_W3p40L3p40_2/w_153_153# a_200_110# 2.41fF
C53 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/w_153_153# a_200_110# 2.41fF
C54 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/a_330_330# a_200_110# 0.65fF
C55 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/w_153_153# a_200_110# 2.41fF
