magic
tech sky130A
timestamp 1616199731
<< nwell >>
rect 200 1464 350 9600
<< mvpmos >>
rect 250 1532 300 9532
<< mvpdiff >>
rect 250 9558 300 9567
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 250 9532 300 9541
rect 250 1523 300 1532
rect 250 1506 258 1523
rect 292 1506 300 1523
rect 250 1497 300 1506
<< mvpdiffc >>
rect 258 9541 292 9558
rect 258 1506 292 1523
<< poly >>
rect 200 1532 250 9532
rect 300 1532 350 9532
<< locali >>
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 250 1506 258 1523
rect 292 1506 300 1523
<< end >>
