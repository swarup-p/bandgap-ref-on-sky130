**.subckt bandgap_ref_cir
XM1 net1 net1 Vrefl GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net2 net1 Vrefr1 GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XQ1 GND GND Vrefl GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ2 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XM10 Vbgp net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XQ3 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ4 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ5 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ6 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ7 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ8 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ9 GND GND Vrefr2 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
R1 Vrefr1 Vrefr2 20k m=1
R2 Vbgp V1 179k m=1
XQ10 GND GND V1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XM3 net2 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
Vdd VDD GND 3.3
XM4 net4 net1 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net3 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
R3 VDD net4 100k m=1
RL Vbgp GND 100Meg m=1
V_en en GND 3.3
XM6 enbar en GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 enbar en VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 net2 en net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM11 net1 enbar GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
**** begin user architecture code


.lib /home/swarup/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt
.include /home/swarup/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130_fd_pr__model__pnp.model.spice
.options savecurrents

*** plot vbgp with variation in supply voltage
.dc vdd 2.7 3.9 0.05
*.control
*run
*plot V(Vbgp)
*.endc

*** plot vbgp with variation in temperature @3.3V
*.dc temp -40 140 1
*.control
*run
*print V(Vbgp)
*plot V(Vbgp)
*.endc

*** plot voltage coefficient
*.dc vdd 2.1 3.6 0.05
*.control
*run
*plot deriv(V(Vbgp))
*.endc

*** plot temperature coefficient
*.dc temp -40 125 1
*.control
*run
*plot deriv(V(Vbgp))/1.2040
*.endc

*** check start up circuit
*Vdd VDD GND PULSE(0 3.3 50us 50us 0us 300us 500us 0)
*.tran 1us 300us
*.control
*run
*plot V(Vdd) V(Vbgp)
*.endc

*** enable pin
*V_en en GND PULSE(0 3.3 0 0 0 10us 20us 0)
*.tran 1u 50us
*.control
*run
*plot V(V_en) V(Vbgp)
*.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.GLOBAL en
.GLOBAL enbar
** flattened .save nodes
.end
