* SPICE3 file created from bgr_a3.ext - technology: sky130A

.lib ../../pre-layout/sky130_fd_pr/models/sky130_tt_bgr.lib.spice tt
.option scale=0.005u
.options savecurrents

X0 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND F sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 C VbiasN VbiasP GND sky130_fd_pr__nfet_g5v0d10v5 w=3000 l=1000
X2 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 G VbiasN VbiasN GND sky130_fd_pr__nfet_g5v0d10v5 w=3000 l=1000
X4 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A  sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X7 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X8 GND I VbiasP GND sky130_fd_pr__nfet_g5v0d10v5 w=600 l=200
X9 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X10 GND VbiasN I GND sky130_fd_pr__nfet_g5v0d10v5 w=600 l=200
X11 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X12 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND A sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X13 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# GND J sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40
X14 VDD VbiasP VbiasN VDD sky130_fd_pr__pfet_g5v0d10v5 w=3000 l=1000
X15 VDD VbiasP VbiasP VDD sky130_fd_pr__pfet_g5v0d10v5 w=3000 l=1000
X16 VDD VbiasP E VDD sky130_fd_pr__pfet_g5v0d10v5 w=3000 l=1000
X17 G en F GND sky130_fd_pr__nfet_g5v0d10v5 w=2400 l=1000
X18 C en B GND sky130_fd_pr__nfet_g5v0d10v5 w=2400 l=1000
X19 Vbgp en E GND sky130_fd_pr__nfet_g5v0d10v5 w=2400 l=1000
X20 A B GND sky130_fd_pr__res_xhigh_po w=70 l=1750
X21 Vbgp H GND sky130_fd_pr__res_xhigh_po w=70 l=8102
X22 VDD I I VDD sky130_fd_pr__pfet_g5v0d10v5 w=100 l=16000
X23 J H GND sky130_fd_pr__res_xhigh_po w=70 l=8102
C0 VbiasN VDD 0.00fF
C1 A J 0.02fF
C2 VbiasN I 1.34fF
C3 C en 0.58fF
C4 G en 0.58fF
C5 VbiasP VDD 1.23fF
C6 A F 0.09fF
C7 VbiasP I 4.85fF
C8 B C 0.06fF
C9 J Vbgp 0.14fF
C10 B Vbgp 0.04fF
C11 E en 0.58fF
C12 A Vbgp 0.89fF
C13 I VDD 0.01fF
C14 E B 0.06fF
C15 VbiasN en 0.23fF
C16 E VDD 0.00fF
C17 VbiasP VbiasN 3.79fF
C18 E C 0.15fF
C19 B en 1.45fF
C20 en GND 16.67fF
C21 VbiasN GND 4.28fF
C22 H GND 0.33fF
C23 Vbgp GND 0.82fF
C24 E GND 0.06fF
C25 B GND 0.89fF
C26 VDD GND 147.24fF
C27 J GND 1.81fF
C28 A GND 3.04fF
C29 F GND 0.10fF

*** plot vbgp with variation in temperature @3.3V
Vdd VDD GND 3.3
V_en en GND 3.3
RLoad Vbgp GND 100Meg
.dc temp -40 140 1
.control
run
print Vbgp
plot V(Vbgp)
.endc
.end
