magic
tech sky130A
timestamp 1615962681
<< nwell >>
rect 0 9600 10000 10000
rect 200 1464 350 9600
rect 700 7630 1336 9600
rect 1486 7630 2122 9600
rect 2272 7630 2908 9600
<< mvnmos >>
rect 768 5779 1268 7279
rect 1554 5779 2054 7279
rect 768 4177 1268 5377
rect 1554 4177 2054 5377
rect 2340 4177 2840 5377
rect 225 1028 325 1328
rect 225 601 325 901
<< mvpmos >>
rect 250 1532 300 9532
rect 768 7749 1268 9249
rect 1554 7749 2054 9249
rect 2340 7749 2840 9249
<< mvndiff >>
rect 733 7222 768 7279
rect 733 7137 742 7222
rect 759 7137 768 7222
rect 733 7037 768 7137
rect 733 6952 742 7037
rect 759 6952 768 7037
rect 733 6852 768 6952
rect 733 6767 742 6852
rect 759 6767 768 6852
rect 733 6667 768 6767
rect 733 6582 742 6667
rect 759 6582 768 6667
rect 733 6482 768 6582
rect 733 6397 742 6482
rect 759 6397 768 6482
rect 733 6297 768 6397
rect 733 6212 742 6297
rect 759 6212 768 6297
rect 733 6112 768 6212
rect 733 6027 742 6112
rect 759 6027 768 6112
rect 733 5927 768 6027
rect 733 5842 742 5927
rect 759 5842 768 5927
rect 733 5779 768 5842
rect 1268 7222 1303 7279
rect 1268 7137 1277 7222
rect 1294 7137 1303 7222
rect 1268 7037 1303 7137
rect 1268 6952 1277 7037
rect 1294 6952 1303 7037
rect 1268 6852 1303 6952
rect 1268 6767 1277 6852
rect 1294 6767 1303 6852
rect 1268 6667 1303 6767
rect 1268 6582 1277 6667
rect 1294 6582 1303 6667
rect 1268 6482 1303 6582
rect 1268 6397 1277 6482
rect 1294 6397 1303 6482
rect 1268 6297 1303 6397
rect 1268 6212 1277 6297
rect 1294 6212 1303 6297
rect 1268 6112 1303 6212
rect 1268 6027 1277 6112
rect 1294 6027 1303 6112
rect 1268 5927 1303 6027
rect 1268 5842 1277 5927
rect 1294 5842 1303 5927
rect 1268 5779 1303 5842
rect 1519 7222 1554 7279
rect 1519 7137 1528 7222
rect 1545 7137 1554 7222
rect 1519 7037 1554 7137
rect 1519 6952 1528 7037
rect 1545 6952 1554 7037
rect 1519 6852 1554 6952
rect 1519 6767 1528 6852
rect 1545 6767 1554 6852
rect 1519 6667 1554 6767
rect 1519 6582 1528 6667
rect 1545 6582 1554 6667
rect 1519 6482 1554 6582
rect 1519 6397 1528 6482
rect 1545 6397 1554 6482
rect 1519 6297 1554 6397
rect 1519 6212 1528 6297
rect 1545 6212 1554 6297
rect 1519 6112 1554 6212
rect 1519 6027 1528 6112
rect 1545 6027 1554 6112
rect 1519 5927 1554 6027
rect 1519 5842 1528 5927
rect 1545 5842 1554 5927
rect 1519 5779 1554 5842
rect 2054 7222 2089 7279
rect 2054 7137 2063 7222
rect 2080 7137 2089 7222
rect 2054 7037 2089 7137
rect 2054 6952 2063 7037
rect 2080 6952 2089 7037
rect 2054 6852 2089 6952
rect 2054 6767 2063 6852
rect 2080 6767 2089 6852
rect 2054 6667 2089 6767
rect 2054 6582 2063 6667
rect 2080 6582 2089 6667
rect 2054 6482 2089 6582
rect 2054 6397 2063 6482
rect 2080 6397 2089 6482
rect 2054 6297 2089 6397
rect 2054 6212 2063 6297
rect 2080 6212 2089 6297
rect 2054 6112 2089 6212
rect 2054 6027 2063 6112
rect 2080 6027 2089 6112
rect 2054 5927 2089 6027
rect 2054 5842 2063 5927
rect 2080 5842 2089 5927
rect 2054 5779 2089 5842
rect 733 5282 768 5377
rect 733 5197 742 5282
rect 759 5197 768 5282
rect 733 5097 768 5197
rect 733 5012 742 5097
rect 759 5012 768 5097
rect 733 4912 768 5012
rect 733 4827 742 4912
rect 759 4827 768 4912
rect 733 4727 768 4827
rect 733 4642 742 4727
rect 759 4642 768 4727
rect 733 4542 768 4642
rect 733 4457 742 4542
rect 759 4457 768 4542
rect 733 4357 768 4457
rect 733 4272 742 4357
rect 759 4272 768 4357
rect 733 4177 768 4272
rect 1268 5282 1303 5377
rect 1268 5197 1277 5282
rect 1294 5197 1303 5282
rect 1268 5097 1303 5197
rect 1268 5012 1277 5097
rect 1294 5012 1303 5097
rect 1268 4912 1303 5012
rect 1268 4827 1277 4912
rect 1294 4827 1303 4912
rect 1268 4727 1303 4827
rect 1268 4642 1277 4727
rect 1294 4642 1303 4727
rect 1268 4542 1303 4642
rect 1268 4457 1277 4542
rect 1294 4457 1303 4542
rect 1268 4357 1303 4457
rect 1268 4272 1277 4357
rect 1294 4272 1303 4357
rect 1268 4177 1303 4272
rect 1519 5282 1554 5377
rect 1519 5197 1528 5282
rect 1545 5197 1554 5282
rect 1519 5097 1554 5197
rect 1519 5012 1528 5097
rect 1545 5012 1554 5097
rect 1519 4912 1554 5012
rect 1519 4827 1528 4912
rect 1545 4827 1554 4912
rect 1519 4727 1554 4827
rect 1519 4642 1528 4727
rect 1545 4642 1554 4727
rect 1519 4542 1554 4642
rect 1519 4457 1528 4542
rect 1545 4457 1554 4542
rect 1519 4357 1554 4457
rect 1519 4272 1528 4357
rect 1545 4272 1554 4357
rect 1519 4177 1554 4272
rect 2054 5282 2089 5377
rect 2054 5197 2063 5282
rect 2080 5197 2089 5282
rect 2054 5097 2089 5197
rect 2054 5012 2063 5097
rect 2080 5012 2089 5097
rect 2054 4912 2089 5012
rect 2054 4827 2063 4912
rect 2080 4827 2089 4912
rect 2054 4727 2089 4827
rect 2054 4642 2063 4727
rect 2080 4642 2089 4727
rect 2054 4542 2089 4642
rect 2054 4457 2063 4542
rect 2080 4457 2089 4542
rect 2054 4357 2089 4457
rect 2054 4272 2063 4357
rect 2080 4272 2089 4357
rect 2054 4177 2089 4272
rect 2305 5282 2340 5377
rect 2305 5197 2314 5282
rect 2331 5197 2340 5282
rect 2305 5097 2340 5197
rect 2305 5012 2314 5097
rect 2331 5012 2340 5097
rect 2305 4912 2340 5012
rect 2305 4827 2314 4912
rect 2331 4827 2340 4912
rect 2305 4727 2340 4827
rect 2305 4642 2314 4727
rect 2331 4642 2340 4727
rect 2305 4542 2340 4642
rect 2305 4457 2314 4542
rect 2331 4457 2340 4542
rect 2305 4357 2340 4457
rect 2305 4272 2314 4357
rect 2331 4272 2340 4357
rect 2305 4177 2340 4272
rect 2840 5282 2875 5377
rect 2840 5197 2849 5282
rect 2866 5197 2875 5282
rect 2840 5097 2875 5197
rect 2840 5012 2849 5097
rect 2866 5012 2875 5097
rect 2840 4912 2875 5012
rect 2840 4827 2849 4912
rect 2866 4827 2875 4912
rect 2840 4727 2875 4827
rect 2840 4642 2849 4727
rect 2866 4642 2875 4727
rect 2840 4542 2875 4642
rect 2840 4457 2849 4542
rect 2866 4457 2875 4542
rect 2840 4357 2875 4457
rect 2840 4272 2849 4357
rect 2866 4272 2875 4357
rect 2840 4177 2875 4272
rect 190 1319 225 1328
rect 190 1228 199 1319
rect 216 1228 225 1319
rect 190 1128 225 1228
rect 190 1037 199 1128
rect 216 1037 225 1128
rect 190 1028 225 1037
rect 325 1319 360 1328
rect 325 1228 334 1319
rect 351 1228 360 1319
rect 325 1128 360 1228
rect 325 1037 334 1128
rect 351 1037 360 1128
rect 325 1028 360 1037
rect 190 892 225 901
rect 190 801 199 892
rect 216 801 225 892
rect 190 701 225 801
rect 190 610 199 701
rect 216 610 225 701
rect 190 601 225 610
rect 325 892 360 901
rect 325 801 334 892
rect 351 801 360 892
rect 325 701 360 801
rect 325 610 334 701
rect 351 610 360 701
rect 325 601 360 610
<< mvpdiff >>
rect 250 9558 300 9567
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 250 9532 300 9541
rect 733 9192 768 9249
rect 733 9107 742 9192
rect 759 9107 768 9192
rect 733 9007 768 9107
rect 733 8922 742 9007
rect 759 8922 768 9007
rect 733 8822 768 8922
rect 733 8737 742 8822
rect 759 8737 768 8822
rect 733 8637 768 8737
rect 733 8552 742 8637
rect 759 8552 768 8637
rect 733 8452 768 8552
rect 733 8367 742 8452
rect 759 8367 768 8452
rect 733 8267 768 8367
rect 733 8182 742 8267
rect 759 8182 768 8267
rect 733 8082 768 8182
rect 733 7997 742 8082
rect 759 7997 768 8082
rect 733 7897 768 7997
rect 733 7812 742 7897
rect 759 7812 768 7897
rect 733 7749 768 7812
rect 1268 9192 1303 9249
rect 1268 9107 1277 9192
rect 1294 9107 1303 9192
rect 1268 9007 1303 9107
rect 1268 8922 1277 9007
rect 1294 8922 1303 9007
rect 1268 8822 1303 8922
rect 1268 8737 1277 8822
rect 1294 8737 1303 8822
rect 1268 8637 1303 8737
rect 1268 8552 1277 8637
rect 1294 8552 1303 8637
rect 1268 8452 1303 8552
rect 1268 8367 1277 8452
rect 1294 8367 1303 8452
rect 1268 8267 1303 8367
rect 1268 8182 1277 8267
rect 1294 8182 1303 8267
rect 1268 8082 1303 8182
rect 1268 7997 1277 8082
rect 1294 7997 1303 8082
rect 1268 7897 1303 7997
rect 1268 7812 1277 7897
rect 1294 7812 1303 7897
rect 1268 7749 1303 7812
rect 1519 9192 1554 9249
rect 1519 9107 1528 9192
rect 1545 9107 1554 9192
rect 1519 9007 1554 9107
rect 1519 8922 1528 9007
rect 1545 8922 1554 9007
rect 1519 8822 1554 8922
rect 1519 8737 1528 8822
rect 1545 8737 1554 8822
rect 1519 8637 1554 8737
rect 1519 8552 1528 8637
rect 1545 8552 1554 8637
rect 1519 8452 1554 8552
rect 1519 8367 1528 8452
rect 1545 8367 1554 8452
rect 1519 8267 1554 8367
rect 1519 8182 1528 8267
rect 1545 8182 1554 8267
rect 1519 8082 1554 8182
rect 1519 7997 1528 8082
rect 1545 7997 1554 8082
rect 1519 7897 1554 7997
rect 1519 7812 1528 7897
rect 1545 7812 1554 7897
rect 1519 7749 1554 7812
rect 2054 9192 2089 9249
rect 2054 9107 2063 9192
rect 2080 9107 2089 9192
rect 2054 9007 2089 9107
rect 2054 8922 2063 9007
rect 2080 8922 2089 9007
rect 2054 8822 2089 8922
rect 2054 8737 2063 8822
rect 2080 8737 2089 8822
rect 2054 8637 2089 8737
rect 2054 8552 2063 8637
rect 2080 8552 2089 8637
rect 2054 8452 2089 8552
rect 2054 8367 2063 8452
rect 2080 8367 2089 8452
rect 2054 8267 2089 8367
rect 2054 8182 2063 8267
rect 2080 8182 2089 8267
rect 2054 8082 2089 8182
rect 2054 7997 2063 8082
rect 2080 7997 2089 8082
rect 2054 7897 2089 7997
rect 2054 7812 2063 7897
rect 2080 7812 2089 7897
rect 2054 7749 2089 7812
rect 2305 9192 2340 9249
rect 2305 9107 2314 9192
rect 2331 9107 2340 9192
rect 2305 9007 2340 9107
rect 2305 8922 2314 9007
rect 2331 8922 2340 9007
rect 2305 8822 2340 8922
rect 2305 8737 2314 8822
rect 2331 8737 2340 8822
rect 2305 8637 2340 8737
rect 2305 8552 2314 8637
rect 2331 8552 2340 8637
rect 2305 8452 2340 8552
rect 2305 8367 2314 8452
rect 2331 8367 2340 8452
rect 2305 8267 2340 8367
rect 2305 8182 2314 8267
rect 2331 8182 2340 8267
rect 2305 8082 2340 8182
rect 2305 7997 2314 8082
rect 2331 7997 2340 8082
rect 2305 7897 2340 7997
rect 2305 7812 2314 7897
rect 2331 7812 2340 7897
rect 2305 7749 2340 7812
rect 2840 9192 2875 9249
rect 2840 9107 2849 9192
rect 2866 9107 2875 9192
rect 2840 9007 2875 9107
rect 2840 8922 2849 9007
rect 2866 8922 2875 9007
rect 2840 8822 2875 8922
rect 2840 8737 2849 8822
rect 2866 8737 2875 8822
rect 2840 8637 2875 8737
rect 2840 8552 2849 8637
rect 2866 8552 2875 8637
rect 2840 8452 2875 8552
rect 2840 8367 2849 8452
rect 2866 8367 2875 8452
rect 2840 8267 2875 8367
rect 2840 8182 2849 8267
rect 2866 8182 2875 8267
rect 2840 8082 2875 8182
rect 2840 7997 2849 8082
rect 2866 7997 2875 8082
rect 2840 7897 2875 7997
rect 2840 7812 2849 7897
rect 2866 7812 2875 7897
rect 2840 7749 2875 7812
rect 250 1523 300 1532
rect 250 1506 258 1523
rect 292 1506 300 1523
rect 250 1497 300 1506
<< mvndiffc >>
rect 742 7137 759 7222
rect 742 6952 759 7037
rect 742 6767 759 6852
rect 742 6582 759 6667
rect 742 6397 759 6482
rect 742 6212 759 6297
rect 742 6027 759 6112
rect 742 5842 759 5927
rect 1277 7137 1294 7222
rect 1277 6952 1294 7037
rect 1277 6767 1294 6852
rect 1277 6582 1294 6667
rect 1277 6397 1294 6482
rect 1277 6212 1294 6297
rect 1277 6027 1294 6112
rect 1277 5842 1294 5927
rect 1528 7137 1545 7222
rect 1528 6952 1545 7037
rect 1528 6767 1545 6852
rect 1528 6582 1545 6667
rect 1528 6397 1545 6482
rect 1528 6212 1545 6297
rect 1528 6027 1545 6112
rect 1528 5842 1545 5927
rect 2063 7137 2080 7222
rect 2063 6952 2080 7037
rect 2063 6767 2080 6852
rect 2063 6582 2080 6667
rect 2063 6397 2080 6482
rect 2063 6212 2080 6297
rect 2063 6027 2080 6112
rect 2063 5842 2080 5927
rect 742 5197 759 5282
rect 742 5012 759 5097
rect 742 4827 759 4912
rect 742 4642 759 4727
rect 742 4457 759 4542
rect 742 4272 759 4357
rect 1277 5197 1294 5282
rect 1277 5012 1294 5097
rect 1277 4827 1294 4912
rect 1277 4642 1294 4727
rect 1277 4457 1294 4542
rect 1277 4272 1294 4357
rect 1528 5197 1545 5282
rect 1528 5012 1545 5097
rect 1528 4827 1545 4912
rect 1528 4642 1545 4727
rect 1528 4457 1545 4542
rect 1528 4272 1545 4357
rect 2063 5197 2080 5282
rect 2063 5012 2080 5097
rect 2063 4827 2080 4912
rect 2063 4642 2080 4727
rect 2063 4457 2080 4542
rect 2063 4272 2080 4357
rect 2314 5197 2331 5282
rect 2314 5012 2331 5097
rect 2314 4827 2331 4912
rect 2314 4642 2331 4727
rect 2314 4457 2331 4542
rect 2314 4272 2331 4357
rect 2849 5197 2866 5282
rect 2849 5012 2866 5097
rect 2849 4827 2866 4912
rect 2849 4642 2866 4727
rect 2849 4457 2866 4542
rect 2849 4272 2866 4357
rect 199 1228 216 1319
rect 199 1037 216 1128
rect 334 1228 351 1319
rect 334 1037 351 1128
rect 199 801 216 892
rect 199 610 216 701
rect 334 801 351 892
rect 334 610 351 701
<< mvpdiffc >>
rect 258 9541 292 9558
rect 742 9107 759 9192
rect 742 8922 759 9007
rect 742 8737 759 8822
rect 742 8552 759 8637
rect 742 8367 759 8452
rect 742 8182 759 8267
rect 742 7997 759 8082
rect 742 7812 759 7897
rect 1277 9107 1294 9192
rect 1277 8922 1294 9007
rect 1277 8737 1294 8822
rect 1277 8552 1294 8637
rect 1277 8367 1294 8452
rect 1277 8182 1294 8267
rect 1277 7997 1294 8082
rect 1277 7812 1294 7897
rect 1528 9107 1545 9192
rect 1528 8922 1545 9007
rect 1528 8737 1545 8822
rect 1528 8552 1545 8637
rect 1528 8367 1545 8452
rect 1528 8182 1545 8267
rect 1528 7997 1545 8082
rect 1528 7812 1545 7897
rect 2063 9107 2080 9192
rect 2063 8922 2080 9007
rect 2063 8737 2080 8822
rect 2063 8552 2080 8637
rect 2063 8367 2080 8452
rect 2063 8182 2080 8267
rect 2063 7997 2080 8082
rect 2063 7812 2080 7897
rect 2314 9107 2331 9192
rect 2314 8922 2331 9007
rect 2314 8737 2331 8822
rect 2314 8552 2331 8637
rect 2314 8367 2331 8452
rect 2314 8182 2331 8267
rect 2314 7997 2331 8082
rect 2314 7812 2331 7897
rect 2849 9107 2866 9192
rect 2849 8922 2866 9007
rect 2849 8737 2866 8822
rect 2849 8552 2866 8637
rect 2849 8367 2866 8452
rect 2849 8182 2866 8267
rect 2849 7997 2866 8082
rect 2849 7812 2866 7897
rect 258 1506 292 1523
<< mvpsubdiff >>
rect 200 300 9800 390
rect 200 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9800 300
rect 200 110 9800 200
<< mvnsubdiff >>
rect 200 9850 9800 9940
rect 200 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9800 9850
rect 200 9660 9800 9750
<< mvpsubdiffcont >>
rect 320 200 420 300
rect 620 200 720 300
rect 920 200 1020 300
rect 1220 200 1320 300
rect 1520 200 1620 300
rect 1820 200 1920 300
rect 2120 200 2220 300
rect 2420 200 2520 300
rect 2720 200 2820 300
rect 3020 200 3120 300
rect 3320 200 3420 300
rect 3620 200 3720 300
rect 3920 200 4020 300
rect 4220 200 4320 300
rect 4520 200 4620 300
rect 4820 200 4920 300
rect 5120 200 5220 300
rect 5420 200 5520 300
rect 5720 200 5820 300
rect 6020 200 6120 300
rect 6320 200 6420 300
rect 6620 200 6720 300
rect 6920 200 7020 300
rect 7220 200 7320 300
rect 7520 200 7620 300
rect 7820 200 7920 300
rect 8120 200 8220 300
rect 8420 200 8520 300
rect 8720 200 8820 300
rect 9020 200 9120 300
rect 9320 200 9420 300
rect 9620 200 9720 300
<< mvnsubdiffcont >>
rect 320 9750 420 9850
rect 620 9750 720 9850
rect 920 9750 1020 9850
rect 1220 9750 1320 9850
rect 1520 9750 1620 9850
rect 1820 9750 1920 9850
rect 2120 9750 2220 9850
rect 2420 9750 2520 9850
rect 2720 9750 2820 9850
rect 3020 9750 3120 9850
rect 3320 9750 3420 9850
rect 3620 9750 3720 9850
rect 3920 9750 4020 9850
rect 4220 9750 4320 9850
rect 4520 9750 4620 9850
rect 4820 9750 4920 9850
rect 5120 9750 5220 9850
rect 5420 9750 5520 9850
rect 5720 9750 5820 9850
rect 6020 9750 6120 9850
rect 6320 9750 6420 9850
rect 6620 9750 6720 9850
rect 6920 9750 7020 9850
rect 7220 9750 7320 9850
rect 7520 9750 7620 9850
rect 7820 9750 7920 9850
rect 8120 9750 8220 9850
rect 8420 9750 8520 9850
rect 8720 9750 8820 9850
rect 9020 9750 9120 9850
rect 9320 9750 9420 9850
rect 9620 9750 9720 9850
<< poly >>
rect 200 1532 250 9532
rect 300 9482 350 9532
rect 300 9382 325 9482
rect 342 9382 350 9482
rect 300 9282 350 9382
rect 300 9182 325 9282
rect 342 9182 350 9282
rect 768 9249 1268 9300
rect 1554 9249 2054 9300
rect 2340 9249 2840 9300
rect 300 9082 350 9182
rect 300 8982 325 9082
rect 342 8982 350 9082
rect 300 8882 350 8982
rect 300 8782 325 8882
rect 342 8782 350 8882
rect 300 8682 350 8782
rect 300 8582 325 8682
rect 342 8582 350 8682
rect 300 8482 350 8582
rect 300 8382 325 8482
rect 342 8382 350 8482
rect 300 8282 350 8382
rect 300 8182 325 8282
rect 342 8182 350 8282
rect 300 8082 350 8182
rect 300 7982 325 8082
rect 342 7982 350 8082
rect 300 7882 350 7982
rect 300 7782 325 7882
rect 342 7782 350 7882
rect 300 7682 350 7782
rect 768 7724 1268 7749
rect 768 7707 828 7724
rect 888 7707 988 7724
rect 1048 7707 1148 7724
rect 1208 7707 1268 7724
rect 768 7698 1268 7707
rect 1554 7724 2054 7749
rect 1554 7707 1614 7724
rect 1674 7707 1774 7724
rect 1834 7707 1934 7724
rect 1994 7707 2054 7724
rect 1554 7698 2054 7707
rect 2340 7724 2840 7749
rect 2340 7707 2400 7724
rect 2460 7707 2560 7724
rect 2620 7707 2720 7724
rect 2780 7707 2840 7724
rect 2340 7698 2840 7707
rect 300 7582 325 7682
rect 342 7582 350 7682
rect 300 7482 350 7582
rect 300 7382 325 7482
rect 342 7382 350 7482
rect 300 7282 350 7382
rect 300 7182 325 7282
rect 342 7182 350 7282
rect 768 7321 1268 7330
rect 768 7304 828 7321
rect 888 7304 988 7321
rect 1048 7304 1148 7321
rect 1208 7304 1268 7321
rect 768 7279 1268 7304
rect 1554 7321 2054 7330
rect 1554 7304 1614 7321
rect 1674 7304 1774 7321
rect 1834 7304 1934 7321
rect 1994 7304 2054 7321
rect 1554 7279 2054 7304
rect 300 7082 350 7182
rect 300 6982 325 7082
rect 342 6982 350 7082
rect 300 6882 350 6982
rect 300 6782 325 6882
rect 342 6782 350 6882
rect 300 6682 350 6782
rect 300 6582 325 6682
rect 342 6582 350 6682
rect 300 6482 350 6582
rect 300 6382 325 6482
rect 342 6382 350 6482
rect 300 6282 350 6382
rect 300 6182 325 6282
rect 342 6182 350 6282
rect 300 6082 350 6182
rect 300 5982 325 6082
rect 342 5982 350 6082
rect 300 5882 350 5982
rect 300 5782 325 5882
rect 342 5782 350 5882
rect 300 5682 350 5782
rect 768 5728 1268 5779
rect 1554 5728 2054 5779
rect 300 5582 325 5682
rect 342 5582 350 5682
rect 300 5482 350 5582
rect 300 5382 325 5482
rect 342 5382 350 5482
rect 300 5282 350 5382
rect 768 5419 1268 5428
rect 768 5402 828 5419
rect 888 5402 988 5419
rect 1048 5402 1148 5419
rect 1208 5402 1268 5419
rect 768 5377 1268 5402
rect 1554 5419 2054 5428
rect 1554 5402 1614 5419
rect 1674 5402 1774 5419
rect 1834 5402 1934 5419
rect 1994 5402 2054 5419
rect 1554 5377 2054 5402
rect 2340 5419 2840 5428
rect 2340 5402 2400 5419
rect 2460 5402 2560 5419
rect 2620 5402 2720 5419
rect 2780 5402 2840 5419
rect 2340 5377 2840 5402
rect 300 5182 325 5282
rect 342 5182 350 5282
rect 300 5082 350 5182
rect 300 4982 325 5082
rect 342 4982 350 5082
rect 300 4882 350 4982
rect 300 4782 325 4882
rect 342 4782 350 4882
rect 300 4682 350 4782
rect 300 4582 325 4682
rect 342 4582 350 4682
rect 300 4482 350 4582
rect 300 4382 325 4482
rect 342 4382 350 4482
rect 300 4282 350 4382
rect 300 4182 325 4282
rect 342 4182 350 4282
rect 300 4082 350 4182
rect 768 4126 1268 4177
rect 1554 4126 2054 4177
rect 2340 4126 2840 4177
rect 300 3982 325 4082
rect 342 3982 350 4082
rect 300 3882 350 3982
rect 300 3782 325 3882
rect 342 3782 350 3882
rect 300 3682 350 3782
rect 300 3582 325 3682
rect 342 3582 350 3682
rect 300 3482 350 3582
rect 300 3382 325 3482
rect 342 3382 350 3482
rect 300 3282 350 3382
rect 300 3182 325 3282
rect 342 3182 350 3282
rect 300 3082 350 3182
rect 300 2982 325 3082
rect 342 2982 350 3082
rect 300 2882 350 2982
rect 300 2782 325 2882
rect 342 2782 350 2882
rect 300 2682 350 2782
rect 300 2582 325 2682
rect 342 2582 350 2682
rect 300 2482 350 2582
rect 300 2382 325 2482
rect 342 2382 350 2482
rect 300 2282 350 2382
rect 300 2182 325 2282
rect 342 2182 350 2282
rect 300 2082 350 2182
rect 300 1982 325 2082
rect 342 1982 350 2082
rect 300 1882 350 1982
rect 300 1782 325 1882
rect 342 1782 350 1882
rect 300 1682 350 1782
rect 300 1582 325 1682
rect 342 1582 350 1682
rect 300 1532 350 1582
rect 225 1370 325 1379
rect 225 1353 235 1370
rect 315 1353 325 1370
rect 225 1328 325 1353
rect 225 977 325 1028
rect 225 901 325 952
rect 225 576 325 601
rect 225 559 235 576
rect 315 559 325 576
rect 225 550 325 559
<< polycont >>
rect 325 9382 342 9482
rect 325 9182 342 9282
rect 325 8982 342 9082
rect 325 8782 342 8882
rect 325 8582 342 8682
rect 325 8382 342 8482
rect 325 8182 342 8282
rect 325 7982 342 8082
rect 325 7782 342 7882
rect 828 7707 888 7724
rect 988 7707 1048 7724
rect 1148 7707 1208 7724
rect 1614 7707 1674 7724
rect 1774 7707 1834 7724
rect 1934 7707 1994 7724
rect 2400 7707 2460 7724
rect 2560 7707 2620 7724
rect 2720 7707 2780 7724
rect 325 7582 342 7682
rect 325 7382 342 7482
rect 325 7182 342 7282
rect 828 7304 888 7321
rect 988 7304 1048 7321
rect 1148 7304 1208 7321
rect 1614 7304 1674 7321
rect 1774 7304 1834 7321
rect 1934 7304 1994 7321
rect 325 6982 342 7082
rect 325 6782 342 6882
rect 325 6582 342 6682
rect 325 6382 342 6482
rect 325 6182 342 6282
rect 325 5982 342 6082
rect 325 5782 342 5882
rect 325 5582 342 5682
rect 325 5382 342 5482
rect 828 5402 888 5419
rect 988 5402 1048 5419
rect 1148 5402 1208 5419
rect 1614 5402 1674 5419
rect 1774 5402 1834 5419
rect 1934 5402 1994 5419
rect 2400 5402 2460 5419
rect 2560 5402 2620 5419
rect 2720 5402 2780 5419
rect 325 5182 342 5282
rect 325 4982 342 5082
rect 325 4782 342 4882
rect 325 4582 342 4682
rect 325 4382 342 4482
rect 325 4182 342 4282
rect 325 3982 342 4082
rect 325 3782 342 3882
rect 325 3582 342 3682
rect 325 3382 342 3482
rect 325 3182 342 3282
rect 325 2982 342 3082
rect 325 2782 342 2882
rect 325 2582 342 2682
rect 325 2382 342 2482
rect 325 2182 342 2282
rect 325 1982 342 2082
rect 325 1782 342 1882
rect 325 1582 342 1682
rect 235 1353 315 1370
rect 235 559 315 576
<< locali >>
rect 100 9850 9900 9940
rect 100 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9900 9850
rect 100 9660 9900 9750
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 325 9482 342 9532
rect 325 9282 342 9382
rect 325 9082 342 9182
rect 325 8882 342 8982
rect 325 8682 342 8782
rect 325 8482 342 8582
rect 325 8282 342 8382
rect 325 8082 342 8182
rect 325 7882 342 7982
rect 325 7682 342 7782
rect 742 9192 759 9660
rect 742 9007 759 9107
rect 742 8822 759 8922
rect 742 8637 759 8737
rect 742 8452 759 8552
rect 742 8267 759 8367
rect 742 8082 759 8182
rect 742 7897 759 7997
rect 742 7749 759 7812
rect 1277 9192 1294 9249
rect 1277 9007 1294 9107
rect 1277 8822 1294 8922
rect 1277 8637 1294 8737
rect 1277 8507 1294 8552
rect 1528 9192 1545 9660
rect 1528 9007 1545 9107
rect 1528 8822 1545 8922
rect 1528 8637 1545 8737
rect 1277 8490 1400 8507
rect 1418 8490 1430 8507
rect 1277 8452 1294 8490
rect 1277 8267 1294 8367
rect 1277 8082 1294 8182
rect 1277 7897 1294 7997
rect 1277 7749 1294 7812
rect 1528 8452 1545 8552
rect 1528 8267 1545 8367
rect 1528 8082 1545 8182
rect 1528 7897 1545 7997
rect 1528 7749 1545 7812
rect 2063 9192 2080 9249
rect 2063 9007 2080 9107
rect 2063 8822 2080 8922
rect 2063 8637 2080 8737
rect 2063 8507 2080 8552
rect 2314 9192 2331 9660
rect 2314 9007 2331 9107
rect 2314 8822 2331 8922
rect 2314 8637 2331 8737
rect 2063 8490 2190 8507
rect 2208 8490 2220 8507
rect 2063 8452 2080 8490
rect 2063 8267 2080 8367
rect 2063 8082 2080 8182
rect 2063 7897 2080 7997
rect 2063 7724 2080 7812
rect 2314 8452 2331 8552
rect 2314 8267 2331 8367
rect 2314 8082 2331 8182
rect 2314 7897 2331 7997
rect 2314 7749 2331 7812
rect 2849 9192 2866 9249
rect 2849 9007 2866 9107
rect 2849 8822 2866 8922
rect 2849 8637 2866 8737
rect 2849 8507 2866 8552
rect 2849 8490 2976 8507
rect 2994 8490 3006 8507
rect 2849 8452 2866 8490
rect 2849 8267 2866 8367
rect 2849 8082 2866 8182
rect 2849 7897 2866 7997
rect 2849 7749 2866 7812
rect 768 7707 828 7724
rect 888 7707 988 7724
rect 1048 7707 1148 7724
rect 1208 7707 1614 7724
rect 1674 7707 1774 7724
rect 1834 7707 1934 7724
rect 1994 7707 2400 7724
rect 2460 7707 2560 7724
rect 2620 7707 2720 7724
rect 2780 7707 2840 7724
rect 325 7482 342 7582
rect 1402 7574 1420 7707
rect 325 7282 342 7382
rect 325 7082 342 7182
rect 325 6882 342 6982
rect 325 6682 342 6782
rect 325 6482 342 6582
rect 325 6282 342 6382
rect 325 6082 342 6182
rect 325 5882 342 5982
rect 325 5682 342 5782
rect 325 5482 342 5582
rect 325 5282 342 5382
rect 325 5082 342 5182
rect 325 4882 342 4982
rect 325 4682 342 4782
rect 325 4482 342 4582
rect 325 4282 342 4382
rect 325 4082 342 4182
rect 325 3882 342 3982
rect 325 3682 342 3782
rect 325 3482 342 3582
rect 325 3282 342 3382
rect 325 3082 342 3182
rect 325 2882 342 2982
rect 325 2682 342 2782
rect 325 2482 342 2582
rect 325 2282 342 2382
rect 325 2082 342 2182
rect 325 1882 342 1982
rect 325 1682 342 1782
rect 325 1523 342 1582
rect 156 1506 258 1523
rect 292 1506 342 1523
rect 390 7557 1420 7574
rect 156 760 173 1506
rect 266 1370 283 1506
rect 225 1353 235 1370
rect 315 1353 325 1370
rect 199 1319 216 1328
rect 199 1128 216 1228
rect 199 973 216 1037
rect 334 1319 351 1328
rect 334 1187 351 1228
rect 390 1187 407 7557
rect 334 1170 407 1187
rect 440 7471 1419 7488
rect 334 1128 351 1170
rect 334 1028 351 1037
rect 199 956 351 973
rect 199 892 216 901
rect 199 760 216 801
rect 156 743 216 760
rect 199 701 216 743
rect 199 601 216 610
rect 334 892 351 956
rect 334 760 351 801
rect 334 743 396 760
rect 414 743 420 760
rect 334 701 351 743
rect 334 601 351 610
rect 440 576 457 7471
rect 1402 7321 1419 7471
rect 768 7304 828 7321
rect 888 7304 988 7321
rect 1048 7304 1148 7321
rect 1208 7304 1614 7321
rect 1674 7304 1774 7321
rect 1834 7304 1934 7321
rect 1994 7304 2054 7321
rect 742 7222 759 7279
rect 742 7037 759 7137
rect 742 6852 759 6952
rect 742 6667 759 6767
rect 742 6482 759 6582
rect 742 6297 759 6397
rect 742 6112 759 6212
rect 742 5927 759 6027
rect 742 5282 759 5842
rect 1277 7222 1294 7304
rect 1277 7037 1294 7137
rect 1277 6852 1294 6952
rect 1277 6667 1294 6767
rect 1277 6537 1294 6582
rect 1528 7222 1545 7279
rect 1528 7037 1545 7137
rect 1528 6852 1545 6952
rect 1528 6667 1545 6767
rect 1277 6520 1400 6537
rect 1418 6520 1430 6537
rect 1277 6482 1294 6520
rect 1277 6297 1294 6397
rect 1277 6112 1294 6212
rect 1277 5927 1294 6027
rect 1277 5779 1294 5842
rect 1528 6482 1545 6582
rect 1528 6297 1545 6397
rect 1528 6112 1545 6212
rect 1528 5927 1545 6027
rect 776 5402 828 5419
rect 888 5402 988 5419
rect 1048 5402 1148 5419
rect 1208 5402 1268 5419
rect 742 5097 759 5197
rect 742 4912 759 5012
rect 742 4727 759 4827
rect 742 4542 759 4642
rect 742 4357 759 4457
rect 742 4177 759 4272
rect 1277 5282 1294 5377
rect 1277 5097 1294 5197
rect 1277 4912 1294 5012
rect 1277 4727 1294 4827
rect 1277 4542 1294 4642
rect 1277 4357 1294 4457
rect 1277 4177 1294 4272
rect 1528 5282 1545 5842
rect 2063 7222 2080 7279
rect 2063 7037 2080 7137
rect 2063 6852 2080 6952
rect 2063 6667 2080 6767
rect 2063 6537 2080 6582
rect 2063 6520 2190 6537
rect 2208 6520 2220 6537
rect 2063 6482 2080 6520
rect 2063 6297 2080 6397
rect 2063 6112 2080 6212
rect 2063 5927 2080 6027
rect 2063 5779 2080 5842
rect 1562 5402 1614 5419
rect 1674 5402 1774 5419
rect 1834 5402 1934 5419
rect 1994 5402 2054 5419
rect 2340 5402 2400 5419
rect 2460 5402 2560 5419
rect 2620 5402 2720 5419
rect 2780 5402 2840 5419
rect 1528 5097 1545 5197
rect 1528 4912 1545 5012
rect 1528 4727 1545 4827
rect 1528 4542 1545 4642
rect 1528 4357 1545 4457
rect 1528 4177 1545 4272
rect 2063 5282 2080 5377
rect 2063 5097 2080 5197
rect 2063 4912 2080 5012
rect 2063 4727 2080 4827
rect 2063 4542 2080 4642
rect 2063 4357 2080 4457
rect 2063 4177 2080 4272
rect 2314 5282 2331 5377
rect 2314 5097 2331 5197
rect 2314 4912 2331 5012
rect 2314 4727 2331 4827
rect 2314 4542 2331 4642
rect 2314 4357 2331 4457
rect 2314 4177 2331 4272
rect 2849 5282 2866 5377
rect 2849 5097 2866 5197
rect 2849 4912 2866 5012
rect 2849 4787 2866 4827
rect 2849 4770 2976 4787
rect 2994 4770 3006 4787
rect 2849 4727 2866 4770
rect 2849 4542 2866 4642
rect 2849 4357 2866 4457
rect 2849 4177 2866 4272
rect 225 559 235 576
rect 315 559 457 576
rect 100 300 9900 390
rect 100 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9900 300
rect 100 110 9900 200
<< viali >>
rect 1400 8490 1418 8507
rect 2190 8490 2208 8507
rect 2976 8490 2994 8507
rect 396 743 414 760
rect 1400 6520 1418 6537
rect 2190 6520 2208 6537
rect 2976 4770 2994 4787
<< metal1 >>
rect 0 9650 10000 9950
rect 1394 8507 1424 8511
rect 1394 8490 1400 8507
rect 1418 8490 1424 8507
rect 1394 6537 1424 8490
rect 1394 6520 1400 6537
rect 1418 6520 1424 6537
rect 1394 6516 1424 6520
rect 2184 8507 2214 8511
rect 2184 8490 2190 8507
rect 2208 8490 2214 8507
rect 2184 6537 2214 8490
rect 2184 6520 2190 6537
rect 2208 6520 2214 6537
rect 2184 6516 2214 6520
rect 2970 8507 3000 8511
rect 2970 8490 2976 8507
rect 2994 8490 3000 8507
rect 2970 4787 3000 8490
rect 2970 4770 2976 4787
rect 2994 4770 3000 4787
rect 2970 4766 3000 4770
rect 1951 2199 1981 2550
rect 2323 1387 2353 2550
rect 2695 2199 2725 2550
rect 3067 1387 3097 2550
rect 3439 2199 3469 2550
rect 3811 1387 3841 2550
rect 4183 2199 4213 2550
rect 4555 1387 4585 2550
rect 2049 1357 2353 1387
rect 2793 1357 3097 1387
rect 3537 1357 3841 1387
rect 4281 1357 4585 1387
rect 390 760 420 764
rect 390 743 396 760
rect 414 743 420 760
rect 390 500 420 743
rect 0 0 10000 500
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8 ~/bandgap-ref-on-sky130/pre-layout/sky130_fd_pr
timestamp 1615375237
transform 1 0 1568 0 1 1718
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 2312 0 1 1718
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 3056 0 1 1718
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 3800 0 1 1718
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 3800 0 1 974
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 3056 0 1 974
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 2312 0 1 974
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 1568 0 1 974
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 674 0 1 2930
box 26 26 770 795
<< end >>
