magic
tech sky130A
timestamp 1616583909
<< mvnmos >>
rect 225 601 325 2101
<< mvndiff >>
rect 190 2060 225 2101
rect 190 1960 199 2060
rect 216 1960 225 2060
rect 190 1940 225 1960
rect 190 1840 199 1940
rect 216 1840 225 1940
rect 190 1820 225 1840
rect 190 1720 199 1820
rect 216 1720 225 1820
rect 190 1700 225 1720
rect 190 1600 199 1700
rect 216 1600 225 1700
rect 190 1580 225 1600
rect 190 1480 199 1580
rect 216 1480 225 1580
rect 190 1460 225 1480
rect 190 1360 199 1460
rect 216 1360 225 1460
rect 190 1340 225 1360
rect 190 1240 199 1340
rect 216 1240 225 1340
rect 190 1220 225 1240
rect 190 1120 199 1220
rect 216 1120 225 1220
rect 190 1100 225 1120
rect 190 1000 199 1100
rect 216 1000 225 1100
rect 190 980 225 1000
rect 190 880 199 980
rect 216 880 225 980
rect 190 860 225 880
rect 190 760 199 860
rect 216 760 225 860
rect 190 740 225 760
rect 190 640 199 740
rect 216 640 225 740
rect 190 601 225 640
rect 325 2060 360 2101
rect 325 1960 334 2060
rect 351 1960 360 2060
rect 325 1940 360 1960
rect 325 1840 334 1940
rect 351 1840 360 1940
rect 325 1820 360 1840
rect 325 1720 334 1820
rect 351 1720 360 1820
rect 325 1700 360 1720
rect 325 1600 334 1700
rect 351 1600 360 1700
rect 325 1580 360 1600
rect 325 1480 334 1580
rect 351 1480 360 1580
rect 325 1460 360 1480
rect 325 1360 334 1460
rect 351 1360 360 1460
rect 325 1340 360 1360
rect 325 1240 334 1340
rect 351 1240 360 1340
rect 325 1220 360 1240
rect 325 1120 334 1220
rect 351 1120 360 1220
rect 325 1100 360 1120
rect 325 1000 334 1100
rect 351 1000 360 1100
rect 325 980 360 1000
rect 325 880 334 980
rect 351 880 360 980
rect 325 860 360 880
rect 325 760 334 860
rect 351 760 360 860
rect 325 740 360 760
rect 325 640 334 740
rect 351 640 360 740
rect 325 601 360 640
<< mvndiffc >>
rect 199 1960 216 2060
rect 199 1840 216 1940
rect 199 1720 216 1820
rect 199 1600 216 1700
rect 199 1480 216 1580
rect 199 1360 216 1460
rect 199 1240 216 1340
rect 199 1120 216 1220
rect 199 1000 216 1100
rect 199 880 216 980
rect 199 760 216 860
rect 199 640 216 740
rect 334 1960 351 2060
rect 334 1840 351 1940
rect 334 1720 351 1820
rect 334 1600 351 1700
rect 334 1480 351 1580
rect 334 1360 351 1460
rect 334 1240 351 1340
rect 334 1120 351 1220
rect 334 1000 351 1100
rect 334 880 351 980
rect 334 760 351 860
rect 334 640 351 740
<< poly >>
rect 225 2101 325 2152
rect 225 550 325 601
<< locali >>
rect 199 2060 216 2101
rect 199 1940 216 1960
rect 199 1820 216 1840
rect 199 1700 216 1720
rect 199 1580 216 1600
rect 199 1460 216 1480
rect 199 1340 216 1360
rect 199 1220 216 1240
rect 199 1100 216 1120
rect 199 980 216 1000
rect 199 860 216 880
rect 199 740 216 760
rect 199 601 216 640
rect 334 2060 351 2101
rect 334 1940 351 1960
rect 334 1820 351 1840
rect 334 1700 351 1720
rect 334 1580 351 1600
rect 334 1460 351 1480
rect 334 1340 351 1360
rect 334 1220 351 1240
rect 334 1100 351 1120
rect 334 980 351 1000
rect 334 860 351 880
rect 334 740 351 760
rect 334 601 351 640
<< end >>
