magic
tech sky130A
timestamp 1616583729
<< mvnmos >>
rect 225 601 725 2101
<< mvndiff >>
rect 190 2060 225 2101
rect 190 1960 199 2060
rect 216 1960 225 2060
rect 190 1940 225 1960
rect 190 1840 199 1940
rect 216 1840 225 1940
rect 190 1820 225 1840
rect 190 1720 199 1820
rect 216 1720 225 1820
rect 190 1700 225 1720
rect 190 1600 199 1700
rect 216 1600 225 1700
rect 190 1580 225 1600
rect 190 1480 199 1580
rect 216 1480 225 1580
rect 190 1460 225 1480
rect 190 1360 199 1460
rect 216 1360 225 1460
rect 190 1340 225 1360
rect 190 1240 199 1340
rect 216 1240 225 1340
rect 190 1220 225 1240
rect 190 1120 199 1220
rect 216 1120 225 1220
rect 190 1100 225 1120
rect 190 1000 199 1100
rect 216 1000 225 1100
rect 190 980 225 1000
rect 190 880 199 980
rect 216 880 225 980
rect 190 860 225 880
rect 190 760 199 860
rect 216 760 225 860
rect 190 740 225 760
rect 190 640 199 740
rect 216 640 225 740
rect 190 601 225 640
rect 725 2060 760 2101
rect 725 1960 734 2060
rect 751 1960 760 2060
rect 725 1940 760 1960
rect 725 1840 734 1940
rect 751 1840 760 1940
rect 725 1820 760 1840
rect 725 1720 734 1820
rect 751 1720 760 1820
rect 725 1700 760 1720
rect 725 1600 734 1700
rect 751 1600 760 1700
rect 725 1580 760 1600
rect 725 1480 734 1580
rect 751 1480 760 1580
rect 725 1460 760 1480
rect 725 1360 734 1460
rect 751 1360 760 1460
rect 725 1340 760 1360
rect 725 1240 734 1340
rect 751 1240 760 1340
rect 725 1220 760 1240
rect 725 1120 734 1220
rect 751 1120 760 1220
rect 725 1100 760 1120
rect 725 1000 734 1100
rect 751 1000 760 1100
rect 725 980 760 1000
rect 725 880 734 980
rect 751 880 760 980
rect 725 860 760 880
rect 725 760 734 860
rect 751 760 760 860
rect 725 740 760 760
rect 725 640 734 740
rect 751 640 760 740
rect 725 601 760 640
<< mvndiffc >>
rect 199 1960 216 2060
rect 199 1840 216 1940
rect 199 1720 216 1820
rect 199 1600 216 1700
rect 199 1480 216 1580
rect 199 1360 216 1460
rect 199 1240 216 1340
rect 199 1120 216 1220
rect 199 1000 216 1100
rect 199 880 216 980
rect 199 760 216 860
rect 199 640 216 740
rect 734 1960 751 2060
rect 734 1840 751 1940
rect 734 1720 751 1820
rect 734 1600 751 1700
rect 734 1480 751 1580
rect 734 1360 751 1460
rect 734 1240 751 1340
rect 734 1120 751 1220
rect 734 1000 751 1100
rect 734 880 751 980
rect 734 760 751 860
rect 734 640 751 740
<< poly >>
rect 225 2101 725 2152
rect 225 550 725 601
<< locali >>
rect 199 2060 216 2101
rect 199 1940 216 1960
rect 199 1820 216 1840
rect 199 1700 216 1720
rect 199 1580 216 1600
rect 199 1460 216 1480
rect 199 1340 216 1360
rect 199 1220 216 1240
rect 199 1100 216 1120
rect 199 980 216 1000
rect 199 860 216 880
rect 199 740 216 760
rect 199 601 216 640
rect 734 2060 751 2101
rect 734 1940 751 1960
rect 734 1820 751 1840
rect 734 1700 751 1720
rect 734 1580 751 1600
rect 734 1460 751 1480
rect 734 1340 751 1360
rect 734 1220 751 1240
rect 734 1100 751 1120
rect 734 980 751 1000
rect 734 860 751 880
rect 734 740 751 760
rect 734 601 751 640
<< end >>
