magic
tech sky130A
timestamp 1615589382
<< nwell >>
rect 0 9600 29104 10000
rect 200 1464 350 9600
<< mvnmos >>
rect 225 1028 325 1328
rect 225 601 325 901
<< mvpmos >>
rect 250 1532 300 9532
<< mvndiff >>
rect 190 1319 225 1328
rect 190 1228 199 1319
rect 216 1228 225 1319
rect 190 1128 225 1228
rect 190 1037 199 1128
rect 216 1037 225 1128
rect 190 1028 225 1037
rect 325 1319 360 1328
rect 325 1228 334 1319
rect 351 1228 360 1319
rect 325 1128 360 1228
rect 325 1037 334 1128
rect 351 1037 360 1128
rect 325 1028 360 1037
rect 190 892 225 901
rect 190 801 199 892
rect 216 801 225 892
rect 190 701 225 801
rect 190 610 199 701
rect 216 610 225 701
rect 190 601 225 610
rect 325 892 360 901
rect 325 801 334 892
rect 351 801 360 892
rect 325 701 360 801
rect 325 610 334 701
rect 351 610 360 701
rect 325 601 360 610
<< mvpdiff >>
rect 250 9558 300 9567
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 250 9532 300 9541
rect 250 1523 300 1532
rect 250 1506 258 1523
rect 292 1506 300 1523
rect 250 1497 300 1506
<< mvndiffc >>
rect 199 1228 216 1319
rect 199 1037 216 1128
rect 334 1228 351 1319
rect 334 1037 351 1128
rect 199 801 216 892
rect 199 610 216 701
rect 334 801 351 892
rect 334 610 351 701
<< mvpdiffc >>
rect 258 9541 292 9558
rect 258 1506 292 1523
<< mvpsubdiff >>
rect 200 300 28904 390
rect 200 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9920 300
rect 10020 200 10220 300
rect 10320 200 10520 300
rect 10620 200 10820 300
rect 10920 200 11120 300
rect 11220 200 11420 300
rect 11520 200 11720 300
rect 11820 200 12020 300
rect 12120 200 12320 300
rect 12420 200 12620 300
rect 12720 200 12920 300
rect 13020 200 13220 300
rect 13320 200 13520 300
rect 13620 200 13820 300
rect 13920 200 14120 300
rect 14220 200 14420 300
rect 14520 200 14720 300
rect 14820 200 15020 300
rect 15120 200 15320 300
rect 15420 200 15620 300
rect 15720 200 15920 300
rect 16020 200 16220 300
rect 16320 200 16520 300
rect 16620 200 16820 300
rect 16920 200 17120 300
rect 17220 200 17420 300
rect 17520 200 17720 300
rect 17820 200 18020 300
rect 18120 200 18320 300
rect 18420 200 18620 300
rect 18720 200 18920 300
rect 19020 200 19220 300
rect 19320 200 19520 300
rect 19620 200 19820 300
rect 19920 200 20120 300
rect 20220 200 20420 300
rect 20520 200 20720 300
rect 20820 200 21020 300
rect 21120 200 21320 300
rect 21420 200 21620 300
rect 21720 200 21920 300
rect 22020 200 22220 300
rect 22320 200 22520 300
rect 22620 200 22820 300
rect 22920 200 23120 300
rect 23220 200 23420 300
rect 23520 200 23720 300
rect 23820 200 24020 300
rect 24120 200 24320 300
rect 24420 200 24620 300
rect 24720 200 24920 300
rect 25020 200 25220 300
rect 25320 200 25520 300
rect 25620 200 25820 300
rect 25920 200 26120 300
rect 26220 200 26420 300
rect 26520 200 26720 300
rect 26820 200 27020 300
rect 27120 200 27320 300
rect 27420 200 27620 300
rect 27720 200 27920 300
rect 28020 200 28220 300
rect 28320 200 28520 300
rect 28620 200 28904 300
rect 200 110 28904 200
<< mvnsubdiff >>
rect 200 9850 28904 9940
rect 200 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9920 9850
rect 10020 9750 10220 9850
rect 10320 9750 10520 9850
rect 10620 9750 10820 9850
rect 10920 9750 11120 9850
rect 11220 9750 11420 9850
rect 11520 9750 11720 9850
rect 11820 9750 12020 9850
rect 12120 9750 12320 9850
rect 12420 9750 12620 9850
rect 12720 9750 12920 9850
rect 13020 9750 13220 9850
rect 13320 9750 13520 9850
rect 13620 9750 13820 9850
rect 13920 9750 14120 9850
rect 14220 9750 14420 9850
rect 14520 9750 14720 9850
rect 14820 9750 15020 9850
rect 15120 9750 15320 9850
rect 15420 9750 15620 9850
rect 15720 9750 15920 9850
rect 16020 9750 16220 9850
rect 16320 9750 16520 9850
rect 16620 9750 16820 9850
rect 16920 9750 17120 9850
rect 17220 9750 17420 9850
rect 17520 9750 17720 9850
rect 17820 9750 18020 9850
rect 18120 9750 18320 9850
rect 18420 9750 18620 9850
rect 18720 9750 18920 9850
rect 19020 9750 19220 9850
rect 19320 9750 19520 9850
rect 19620 9750 19820 9850
rect 19920 9750 20120 9850
rect 20220 9750 20420 9850
rect 20520 9750 20720 9850
rect 20820 9750 21020 9850
rect 21120 9750 21320 9850
rect 21420 9750 21620 9850
rect 21720 9750 21920 9850
rect 22020 9750 22220 9850
rect 22320 9750 22520 9850
rect 22620 9750 22820 9850
rect 22920 9750 23120 9850
rect 23220 9750 23420 9850
rect 23520 9750 23720 9850
rect 23820 9750 24020 9850
rect 24120 9750 24320 9850
rect 24420 9750 24620 9850
rect 24720 9750 24920 9850
rect 25020 9750 25220 9850
rect 25320 9750 25520 9850
rect 25620 9750 25820 9850
rect 25920 9750 26120 9850
rect 26220 9750 26420 9850
rect 26520 9750 26720 9850
rect 26820 9750 27020 9850
rect 27120 9750 27320 9850
rect 27420 9750 27620 9850
rect 27720 9750 27920 9850
rect 28020 9750 28220 9850
rect 28320 9750 28520 9850
rect 28620 9750 28904 9850
rect 200 9660 28904 9750
<< mvpsubdiffcont >>
rect 320 200 420 300
rect 620 200 720 300
rect 920 200 1020 300
rect 1220 200 1320 300
rect 1520 200 1620 300
rect 1820 200 1920 300
rect 2120 200 2220 300
rect 2420 200 2520 300
rect 2720 200 2820 300
rect 3020 200 3120 300
rect 3320 200 3420 300
rect 3620 200 3720 300
rect 3920 200 4020 300
rect 4220 200 4320 300
rect 4520 200 4620 300
rect 4820 200 4920 300
rect 5120 200 5220 300
rect 5420 200 5520 300
rect 5720 200 5820 300
rect 6020 200 6120 300
rect 6320 200 6420 300
rect 6620 200 6720 300
rect 6920 200 7020 300
rect 7220 200 7320 300
rect 7520 200 7620 300
rect 7820 200 7920 300
rect 8120 200 8220 300
rect 8420 200 8520 300
rect 8720 200 8820 300
rect 9020 200 9120 300
rect 9320 200 9420 300
rect 9620 200 9720 300
rect 9920 200 10020 300
rect 10220 200 10320 300
rect 10520 200 10620 300
rect 10820 200 10920 300
rect 11120 200 11220 300
rect 11420 200 11520 300
rect 11720 200 11820 300
rect 12020 200 12120 300
rect 12320 200 12420 300
rect 12620 200 12720 300
rect 12920 200 13020 300
rect 13220 200 13320 300
rect 13520 200 13620 300
rect 13820 200 13920 300
rect 14120 200 14220 300
rect 14420 200 14520 300
rect 14720 200 14820 300
rect 15020 200 15120 300
rect 15320 200 15420 300
rect 15620 200 15720 300
rect 15920 200 16020 300
rect 16220 200 16320 300
rect 16520 200 16620 300
rect 16820 200 16920 300
rect 17120 200 17220 300
rect 17420 200 17520 300
rect 17720 200 17820 300
rect 18020 200 18120 300
rect 18320 200 18420 300
rect 18620 200 18720 300
rect 18920 200 19020 300
rect 19220 200 19320 300
rect 19520 200 19620 300
rect 19820 200 19920 300
rect 20120 200 20220 300
rect 20420 200 20520 300
rect 20720 200 20820 300
rect 21020 200 21120 300
rect 21320 200 21420 300
rect 21620 200 21720 300
rect 21920 200 22020 300
rect 22220 200 22320 300
rect 22520 200 22620 300
rect 22820 200 22920 300
rect 23120 200 23220 300
rect 23420 200 23520 300
rect 23720 200 23820 300
rect 24020 200 24120 300
rect 24320 200 24420 300
rect 24620 200 24720 300
rect 24920 200 25020 300
rect 25220 200 25320 300
rect 25520 200 25620 300
rect 25820 200 25920 300
rect 26120 200 26220 300
rect 26420 200 26520 300
rect 26720 200 26820 300
rect 27020 200 27120 300
rect 27320 200 27420 300
rect 27620 200 27720 300
rect 27920 200 28020 300
rect 28220 200 28320 300
rect 28520 200 28620 300
<< mvnsubdiffcont >>
rect 320 9750 420 9850
rect 620 9750 720 9850
rect 920 9750 1020 9850
rect 1220 9750 1320 9850
rect 1520 9750 1620 9850
rect 1820 9750 1920 9850
rect 2120 9750 2220 9850
rect 2420 9750 2520 9850
rect 2720 9750 2820 9850
rect 3020 9750 3120 9850
rect 3320 9750 3420 9850
rect 3620 9750 3720 9850
rect 3920 9750 4020 9850
rect 4220 9750 4320 9850
rect 4520 9750 4620 9850
rect 4820 9750 4920 9850
rect 5120 9750 5220 9850
rect 5420 9750 5520 9850
rect 5720 9750 5820 9850
rect 6020 9750 6120 9850
rect 6320 9750 6420 9850
rect 6620 9750 6720 9850
rect 6920 9750 7020 9850
rect 7220 9750 7320 9850
rect 7520 9750 7620 9850
rect 7820 9750 7920 9850
rect 8120 9750 8220 9850
rect 8420 9750 8520 9850
rect 8720 9750 8820 9850
rect 9020 9750 9120 9850
rect 9320 9750 9420 9850
rect 9620 9750 9720 9850
rect 9920 9750 10020 9850
rect 10220 9750 10320 9850
rect 10520 9750 10620 9850
rect 10820 9750 10920 9850
rect 11120 9750 11220 9850
rect 11420 9750 11520 9850
rect 11720 9750 11820 9850
rect 12020 9750 12120 9850
rect 12320 9750 12420 9850
rect 12620 9750 12720 9850
rect 12920 9750 13020 9850
rect 13220 9750 13320 9850
rect 13520 9750 13620 9850
rect 13820 9750 13920 9850
rect 14120 9750 14220 9850
rect 14420 9750 14520 9850
rect 14720 9750 14820 9850
rect 15020 9750 15120 9850
rect 15320 9750 15420 9850
rect 15620 9750 15720 9850
rect 15920 9750 16020 9850
rect 16220 9750 16320 9850
rect 16520 9750 16620 9850
rect 16820 9750 16920 9850
rect 17120 9750 17220 9850
rect 17420 9750 17520 9850
rect 17720 9750 17820 9850
rect 18020 9750 18120 9850
rect 18320 9750 18420 9850
rect 18620 9750 18720 9850
rect 18920 9750 19020 9850
rect 19220 9750 19320 9850
rect 19520 9750 19620 9850
rect 19820 9750 19920 9850
rect 20120 9750 20220 9850
rect 20420 9750 20520 9850
rect 20720 9750 20820 9850
rect 21020 9750 21120 9850
rect 21320 9750 21420 9850
rect 21620 9750 21720 9850
rect 21920 9750 22020 9850
rect 22220 9750 22320 9850
rect 22520 9750 22620 9850
rect 22820 9750 22920 9850
rect 23120 9750 23220 9850
rect 23420 9750 23520 9850
rect 23720 9750 23820 9850
rect 24020 9750 24120 9850
rect 24320 9750 24420 9850
rect 24620 9750 24720 9850
rect 24920 9750 25020 9850
rect 25220 9750 25320 9850
rect 25520 9750 25620 9850
rect 25820 9750 25920 9850
rect 26120 9750 26220 9850
rect 26420 9750 26520 9850
rect 26720 9750 26820 9850
rect 27020 9750 27120 9850
rect 27320 9750 27420 9850
rect 27620 9750 27720 9850
rect 27920 9750 28020 9850
rect 28220 9750 28320 9850
rect 28520 9750 28620 9850
<< poly >>
rect 200 1532 250 9532
rect 300 5566 350 9532
rect 300 5532 325 5566
rect 342 5532 350 5566
rect 300 1532 350 5532
rect 225 1370 325 1379
rect 225 1353 258 1370
rect 292 1353 325 1370
rect 225 1328 325 1353
rect 225 977 325 1028
rect 225 901 325 952
rect 225 576 325 601
rect 225 559 258 576
rect 292 559 325 576
rect 225 550 325 559
<< polycont >>
rect 325 5532 342 5566
rect 258 1353 292 1370
rect 258 559 292 576
<< locali >>
rect 100 9850 29004 9940
rect 100 9750 320 9850
rect 420 9750 620 9850
rect 720 9750 920 9850
rect 1020 9750 1220 9850
rect 1320 9750 1520 9850
rect 1620 9750 1820 9850
rect 1920 9750 2120 9850
rect 2220 9750 2420 9850
rect 2520 9750 2720 9850
rect 2820 9750 3020 9850
rect 3120 9750 3320 9850
rect 3420 9750 3620 9850
rect 3720 9750 3920 9850
rect 4020 9750 4220 9850
rect 4320 9750 4520 9850
rect 4620 9750 4820 9850
rect 4920 9750 5120 9850
rect 5220 9750 5420 9850
rect 5520 9750 5720 9850
rect 5820 9750 6020 9850
rect 6120 9750 6320 9850
rect 6420 9750 6620 9850
rect 6720 9750 6920 9850
rect 7020 9750 7220 9850
rect 7320 9750 7520 9850
rect 7620 9750 7820 9850
rect 7920 9750 8120 9850
rect 8220 9750 8420 9850
rect 8520 9750 8720 9850
rect 8820 9750 9020 9850
rect 9120 9750 9320 9850
rect 9420 9750 9620 9850
rect 9720 9750 9920 9850
rect 10020 9750 10220 9850
rect 10320 9750 10520 9850
rect 10620 9750 10820 9850
rect 10920 9750 11120 9850
rect 11220 9750 11420 9850
rect 11520 9750 11720 9850
rect 11820 9750 12020 9850
rect 12120 9750 12320 9850
rect 12420 9750 12620 9850
rect 12720 9750 12920 9850
rect 13020 9750 13220 9850
rect 13320 9750 13520 9850
rect 13620 9750 13820 9850
rect 13920 9750 14120 9850
rect 14220 9750 14420 9850
rect 14520 9750 14720 9850
rect 14820 9750 15020 9850
rect 15120 9750 15320 9850
rect 15420 9750 15620 9850
rect 15720 9750 15920 9850
rect 16020 9750 16220 9850
rect 16320 9750 16520 9850
rect 16620 9750 16820 9850
rect 16920 9750 17120 9850
rect 17220 9750 17420 9850
rect 17520 9750 17720 9850
rect 17820 9750 18020 9850
rect 18120 9750 18320 9850
rect 18420 9750 18620 9850
rect 18720 9750 18920 9850
rect 19020 9750 19220 9850
rect 19320 9750 19520 9850
rect 19620 9750 19820 9850
rect 19920 9750 20120 9850
rect 20220 9750 20420 9850
rect 20520 9750 20720 9850
rect 20820 9750 21020 9850
rect 21120 9750 21320 9850
rect 21420 9750 21620 9850
rect 21720 9750 21920 9850
rect 22020 9750 22220 9850
rect 22320 9750 22520 9850
rect 22620 9750 22820 9850
rect 22920 9750 23120 9850
rect 23220 9750 23420 9850
rect 23520 9750 23720 9850
rect 23820 9750 24020 9850
rect 24120 9750 24320 9850
rect 24420 9750 24620 9850
rect 24720 9750 24920 9850
rect 25020 9750 25220 9850
rect 25320 9750 25520 9850
rect 25620 9750 25820 9850
rect 25920 9750 26120 9850
rect 26220 9750 26420 9850
rect 26520 9750 26720 9850
rect 26820 9750 27020 9850
rect 27120 9750 27320 9850
rect 27420 9750 27620 9850
rect 27720 9750 27920 9850
rect 28020 9750 28220 9850
rect 28320 9750 28520 9850
rect 28620 9750 29004 9850
rect 100 9660 29004 9750
rect 258 9558 292 9660
rect 250 9541 258 9558
rect 292 9541 300 9558
rect 325 5566 342 5584
rect 325 1523 342 5532
rect 250 1506 258 1523
rect 292 1506 342 1523
rect 267 1370 284 1506
rect 163 1353 258 1370
rect 292 1353 301 1370
rect 163 761 180 1353
rect 199 1319 216 1328
rect 199 1128 216 1228
rect 199 973 216 1037
rect 334 1319 351 1328
rect 334 1187 351 1228
rect 334 1170 400 1187
rect 334 1128 351 1170
rect 334 1028 351 1037
rect 199 956 351 973
rect 199 892 216 901
rect 199 761 216 801
rect 163 744 216 761
rect 199 701 216 744
rect 199 601 216 610
rect 334 892 351 956
rect 334 761 351 801
rect 334 744 406 761
rect 424 744 430 761
rect 334 701 351 744
rect 334 601 351 610
rect 249 559 258 576
rect 292 559 455 576
rect 100 300 29004 390
rect 100 200 320 300
rect 420 200 620 300
rect 720 200 920 300
rect 1020 200 1220 300
rect 1320 200 1520 300
rect 1620 200 1820 300
rect 1920 200 2120 300
rect 2220 200 2420 300
rect 2520 200 2720 300
rect 2820 200 3020 300
rect 3120 200 3320 300
rect 3420 200 3620 300
rect 3720 200 3920 300
rect 4020 200 4220 300
rect 4320 200 4520 300
rect 4620 200 4820 300
rect 4920 200 5120 300
rect 5220 200 5420 300
rect 5520 200 5720 300
rect 5820 200 6020 300
rect 6120 200 6320 300
rect 6420 200 6620 300
rect 6720 200 6920 300
rect 7020 200 7220 300
rect 7320 200 7520 300
rect 7620 200 7820 300
rect 7920 200 8120 300
rect 8220 200 8420 300
rect 8520 200 8720 300
rect 8820 200 9020 300
rect 9120 200 9320 300
rect 9420 200 9620 300
rect 9720 200 9920 300
rect 10020 200 10220 300
rect 10320 200 10520 300
rect 10620 200 10820 300
rect 10920 200 11120 300
rect 11220 200 11420 300
rect 11520 200 11720 300
rect 11820 200 12020 300
rect 12120 200 12320 300
rect 12420 200 12620 300
rect 12720 200 12920 300
rect 13020 200 13220 300
rect 13320 200 13520 300
rect 13620 200 13820 300
rect 13920 200 14120 300
rect 14220 200 14420 300
rect 14520 200 14720 300
rect 14820 200 15020 300
rect 15120 200 15320 300
rect 15420 200 15620 300
rect 15720 200 15920 300
rect 16020 200 16220 300
rect 16320 200 16520 300
rect 16620 200 16820 300
rect 16920 200 17120 300
rect 17220 200 17420 300
rect 17520 200 17720 300
rect 17820 200 18020 300
rect 18120 200 18320 300
rect 18420 200 18620 300
rect 18720 200 18920 300
rect 19020 200 19220 300
rect 19320 200 19520 300
rect 19620 200 19820 300
rect 19920 200 20120 300
rect 20220 200 20420 300
rect 20520 200 20720 300
rect 20820 200 21020 300
rect 21120 200 21320 300
rect 21420 200 21620 300
rect 21720 200 21920 300
rect 22020 200 22220 300
rect 22320 200 22520 300
rect 22620 200 22820 300
rect 22920 200 23120 300
rect 23220 200 23420 300
rect 23520 200 23720 300
rect 23820 200 24020 300
rect 24120 200 24320 300
rect 24420 200 24620 300
rect 24720 200 24920 300
rect 25020 200 25220 300
rect 25320 200 25520 300
rect 25620 200 25820 300
rect 25920 200 26120 300
rect 26220 200 26420 300
rect 26520 200 26720 300
rect 26820 200 27020 300
rect 27120 200 27320 300
rect 27420 200 27620 300
rect 27720 200 27920 300
rect 28020 200 28220 300
rect 28320 200 28520 300
rect 28620 200 29004 300
rect 100 110 29004 200
<< viali >>
rect 406 744 424 761
<< metal1 >>
rect 0 9650 29104 9950
rect 400 761 430 764
rect 400 744 406 761
rect 424 744 430 761
rect 400 500 430 744
rect 0 0 29104 500
<< labels >>
rlabel locali 445 568 445 568 1 VbiasN
rlabel locali 390 1178 390 1178 1 VbiasP
<< end >>
