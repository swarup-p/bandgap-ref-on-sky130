magic
tech sky130A
timestamp 1616538694
<< mvnmos >>
rect 225 601 825 5101
<< mvndiff >>
rect 190 5060 225 5101
rect 190 4960 199 5060
rect 216 4960 225 5060
rect 190 4940 225 4960
rect 190 4840 199 4940
rect 216 4840 225 4940
rect 190 4820 225 4840
rect 190 4720 199 4820
rect 216 4720 225 4820
rect 190 4700 225 4720
rect 190 4600 199 4700
rect 216 4600 225 4700
rect 190 4580 225 4600
rect 190 4480 199 4580
rect 216 4480 225 4580
rect 190 4460 225 4480
rect 190 4360 199 4460
rect 216 4360 225 4460
rect 190 4340 225 4360
rect 190 4240 199 4340
rect 216 4240 225 4340
rect 190 4220 225 4240
rect 190 4120 199 4220
rect 216 4120 225 4220
rect 190 4100 225 4120
rect 190 4000 199 4100
rect 216 4000 225 4100
rect 190 3980 225 4000
rect 190 3880 199 3980
rect 216 3880 225 3980
rect 190 3860 225 3880
rect 190 3760 199 3860
rect 216 3760 225 3860
rect 190 3740 225 3760
rect 190 3640 199 3740
rect 216 3640 225 3740
rect 190 3620 225 3640
rect 190 3520 199 3620
rect 216 3520 225 3620
rect 190 3500 225 3520
rect 190 3400 199 3500
rect 216 3400 225 3500
rect 190 3380 225 3400
rect 190 3280 199 3380
rect 216 3280 225 3380
rect 190 3260 225 3280
rect 190 3160 199 3260
rect 216 3160 225 3260
rect 190 3140 225 3160
rect 190 3040 199 3140
rect 216 3040 225 3140
rect 190 3020 225 3040
rect 190 2920 199 3020
rect 216 2920 225 3020
rect 190 2900 225 2920
rect 190 2800 199 2900
rect 216 2800 225 2900
rect 190 2780 225 2800
rect 190 2680 199 2780
rect 216 2680 225 2780
rect 190 2660 225 2680
rect 190 2560 199 2660
rect 216 2560 225 2660
rect 190 2540 225 2560
rect 190 2440 199 2540
rect 216 2440 225 2540
rect 190 2420 225 2440
rect 190 2320 199 2420
rect 216 2320 225 2420
rect 190 2300 225 2320
rect 190 2200 199 2300
rect 216 2200 225 2300
rect 190 2180 225 2200
rect 190 2080 199 2180
rect 216 2080 225 2180
rect 190 2060 225 2080
rect 190 1960 199 2060
rect 216 1960 225 2060
rect 190 1940 225 1960
rect 190 1840 199 1940
rect 216 1840 225 1940
rect 190 1820 225 1840
rect 190 1720 199 1820
rect 216 1720 225 1820
rect 190 1700 225 1720
rect 190 1600 199 1700
rect 216 1600 225 1700
rect 190 1580 225 1600
rect 190 1480 199 1580
rect 216 1480 225 1580
rect 190 1460 225 1480
rect 190 1360 199 1460
rect 216 1360 225 1460
rect 190 1340 225 1360
rect 190 1240 199 1340
rect 216 1240 225 1340
rect 190 1220 225 1240
rect 190 1120 199 1220
rect 216 1120 225 1220
rect 190 1100 225 1120
rect 190 1000 199 1100
rect 216 1000 225 1100
rect 190 980 225 1000
rect 190 880 199 980
rect 216 880 225 980
rect 190 860 225 880
rect 190 760 199 860
rect 216 760 225 860
rect 190 740 225 760
rect 190 640 199 740
rect 216 640 225 740
rect 190 601 225 640
rect 825 5060 860 5101
rect 825 4960 834 5060
rect 851 4960 860 5060
rect 825 4940 860 4960
rect 825 4840 834 4940
rect 851 4840 860 4940
rect 825 4820 860 4840
rect 825 4720 834 4820
rect 851 4720 860 4820
rect 825 4700 860 4720
rect 825 4600 834 4700
rect 851 4600 860 4700
rect 825 4580 860 4600
rect 825 4480 834 4580
rect 851 4480 860 4580
rect 825 4460 860 4480
rect 825 4360 834 4460
rect 851 4360 860 4460
rect 825 4340 860 4360
rect 825 4240 834 4340
rect 851 4240 860 4340
rect 825 4220 860 4240
rect 825 4120 834 4220
rect 851 4120 860 4220
rect 825 4100 860 4120
rect 825 4000 834 4100
rect 851 4000 860 4100
rect 825 3980 860 4000
rect 825 3880 834 3980
rect 851 3880 860 3980
rect 825 3860 860 3880
rect 825 3760 834 3860
rect 851 3760 860 3860
rect 825 3740 860 3760
rect 825 3640 834 3740
rect 851 3640 860 3740
rect 825 3620 860 3640
rect 825 3520 834 3620
rect 851 3520 860 3620
rect 825 3500 860 3520
rect 825 3400 834 3500
rect 851 3400 860 3500
rect 825 3380 860 3400
rect 825 3280 834 3380
rect 851 3280 860 3380
rect 825 3260 860 3280
rect 825 3160 834 3260
rect 851 3160 860 3260
rect 825 3140 860 3160
rect 825 3040 834 3140
rect 851 3040 860 3140
rect 825 3020 860 3040
rect 825 2920 834 3020
rect 851 2920 860 3020
rect 825 2900 860 2920
rect 825 2800 834 2900
rect 851 2800 860 2900
rect 825 2780 860 2800
rect 825 2680 834 2780
rect 851 2680 860 2780
rect 825 2660 860 2680
rect 825 2560 834 2660
rect 851 2560 860 2660
rect 825 2540 860 2560
rect 825 2440 834 2540
rect 851 2440 860 2540
rect 825 2420 860 2440
rect 825 2320 834 2420
rect 851 2320 860 2420
rect 825 2300 860 2320
rect 825 2200 834 2300
rect 851 2200 860 2300
rect 825 2180 860 2200
rect 825 2080 834 2180
rect 851 2080 860 2180
rect 825 2060 860 2080
rect 825 1960 834 2060
rect 851 1960 860 2060
rect 825 1940 860 1960
rect 825 1840 834 1940
rect 851 1840 860 1940
rect 825 1820 860 1840
rect 825 1720 834 1820
rect 851 1720 860 1820
rect 825 1700 860 1720
rect 825 1600 834 1700
rect 851 1600 860 1700
rect 825 1580 860 1600
rect 825 1480 834 1580
rect 851 1480 860 1580
rect 825 1460 860 1480
rect 825 1360 834 1460
rect 851 1360 860 1460
rect 825 1340 860 1360
rect 825 1240 834 1340
rect 851 1240 860 1340
rect 825 1220 860 1240
rect 825 1120 834 1220
rect 851 1120 860 1220
rect 825 1100 860 1120
rect 825 1000 834 1100
rect 851 1000 860 1100
rect 825 980 860 1000
rect 825 880 834 980
rect 851 880 860 980
rect 825 860 860 880
rect 825 760 834 860
rect 851 760 860 860
rect 825 740 860 760
rect 825 640 834 740
rect 851 640 860 740
rect 825 601 860 640
<< mvndiffc >>
rect 199 4960 216 5060
rect 199 4840 216 4940
rect 199 4720 216 4820
rect 199 4600 216 4700
rect 199 4480 216 4580
rect 199 4360 216 4460
rect 199 4240 216 4340
rect 199 4120 216 4220
rect 199 4000 216 4100
rect 199 3880 216 3980
rect 199 3760 216 3860
rect 199 3640 216 3740
rect 199 3520 216 3620
rect 199 3400 216 3500
rect 199 3280 216 3380
rect 199 3160 216 3260
rect 199 3040 216 3140
rect 199 2920 216 3020
rect 199 2800 216 2900
rect 199 2680 216 2780
rect 199 2560 216 2660
rect 199 2440 216 2540
rect 199 2320 216 2420
rect 199 2200 216 2300
rect 199 2080 216 2180
rect 199 1960 216 2060
rect 199 1840 216 1940
rect 199 1720 216 1820
rect 199 1600 216 1700
rect 199 1480 216 1580
rect 199 1360 216 1460
rect 199 1240 216 1340
rect 199 1120 216 1220
rect 199 1000 216 1100
rect 199 880 216 980
rect 199 760 216 860
rect 199 640 216 740
rect 834 4960 851 5060
rect 834 4840 851 4940
rect 834 4720 851 4820
rect 834 4600 851 4700
rect 834 4480 851 4580
rect 834 4360 851 4460
rect 834 4240 851 4340
rect 834 4120 851 4220
rect 834 4000 851 4100
rect 834 3880 851 3980
rect 834 3760 851 3860
rect 834 3640 851 3740
rect 834 3520 851 3620
rect 834 3400 851 3500
rect 834 3280 851 3380
rect 834 3160 851 3260
rect 834 3040 851 3140
rect 834 2920 851 3020
rect 834 2800 851 2900
rect 834 2680 851 2780
rect 834 2560 851 2660
rect 834 2440 851 2540
rect 834 2320 851 2420
rect 834 2200 851 2300
rect 834 2080 851 2180
rect 834 1960 851 2060
rect 834 1840 851 1940
rect 834 1720 851 1820
rect 834 1600 851 1700
rect 834 1480 851 1580
rect 834 1360 851 1460
rect 834 1240 851 1340
rect 834 1120 851 1220
rect 834 1000 851 1100
rect 834 880 851 980
rect 834 760 851 860
rect 834 640 851 740
<< poly >>
rect 225 5101 825 5152
rect 225 550 825 601
<< locali >>
rect 199 5060 216 5101
rect 199 4940 216 4960
rect 199 4820 216 4840
rect 199 4700 216 4720
rect 199 4580 216 4600
rect 199 4460 216 4480
rect 199 4340 216 4360
rect 199 4220 216 4240
rect 199 4100 216 4120
rect 199 3980 216 4000
rect 199 3860 216 3880
rect 199 3740 216 3760
rect 199 3620 216 3640
rect 199 3500 216 3520
rect 199 3380 216 3400
rect 199 3260 216 3280
rect 199 3140 216 3160
rect 199 3020 216 3040
rect 199 2900 216 2920
rect 199 2780 216 2800
rect 199 2660 216 2680
rect 199 2540 216 2560
rect 199 2420 216 2440
rect 199 2300 216 2320
rect 199 2180 216 2200
rect 199 2060 216 2080
rect 199 1940 216 1960
rect 199 1820 216 1840
rect 199 1700 216 1720
rect 199 1580 216 1600
rect 199 1460 216 1480
rect 199 1340 216 1360
rect 199 1220 216 1240
rect 199 1100 216 1120
rect 199 980 216 1000
rect 199 860 216 880
rect 199 740 216 760
rect 199 601 216 640
rect 834 5060 851 5101
rect 834 4940 851 4960
rect 834 4820 851 4840
rect 834 4700 851 4720
rect 834 4580 851 4600
rect 834 4460 851 4480
rect 834 4340 851 4360
rect 834 4220 851 4240
rect 834 4100 851 4120
rect 834 3980 851 4000
rect 834 3860 851 3880
rect 834 3740 851 3760
rect 834 3620 851 3640
rect 834 3500 851 3520
rect 834 3380 851 3400
rect 834 3260 851 3280
rect 834 3140 851 3160
rect 834 3020 851 3040
rect 834 2900 851 2920
rect 834 2780 851 2800
rect 834 2660 851 2680
rect 834 2540 851 2560
rect 834 2420 851 2440
rect 834 2300 851 2320
rect 834 2180 851 2200
rect 834 2060 851 2080
rect 834 1940 851 1960
rect 834 1820 851 1840
rect 834 1700 851 1720
rect 834 1580 851 1600
rect 834 1460 851 1480
rect 834 1340 851 1360
rect 834 1220 851 1240
rect 834 1100 851 1120
rect 834 980 851 1000
rect 834 860 851 880
rect 834 740 851 760
rect 834 601 851 640
<< end >>
