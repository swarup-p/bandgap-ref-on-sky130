magic
tech sky130A
timestamp 1616028282
<< xpolycontact >>
rect 0 1431 216 1466
rect 1026 1431 1242 1466
rect 0 1272 216 1307
rect 1026 1272 1242 1307
rect 0 1113 216 1148
rect 1026 1113 1242 1148
rect 2700 1026 2735 1242
rect 0 954 216 989
rect 1026 954 1242 989
rect 0 795 216 830
rect 1026 795 1242 830
rect 0 636 216 671
rect 1026 636 1242 671
rect 0 477 216 512
rect 1026 477 1242 512
rect 0 318 216 353
rect 1026 318 1242 353
rect 0 159 216 194
rect 1026 159 1242 194
rect 0 0 216 35
rect 1026 0 1242 35
rect 2700 0 2735 216
rect 2859 1026 2894 1242
rect 2859 0 2894 216
rect 3018 1026 3053 1242
rect 3018 0 3053 216
rect 3177 1026 3212 1242
rect 3177 0 3212 216
rect 3336 1026 3371 1242
rect 3336 0 3371 216
rect 3495 1026 3530 1242
rect 3495 0 3530 216
rect 3654 1026 3689 1242
rect 3654 0 3689 216
rect 3813 1026 3848 1242
rect 3813 0 3848 216
rect 3972 1026 4007 1242
rect 3972 0 4007 216
rect 4131 1026 4166 1242
rect 4131 0 4166 216
<< xpolyres >>
rect 216 1431 1026 1466
rect 216 1272 1026 1307
rect 216 1113 1026 1148
rect 216 954 1026 989
rect 216 795 1026 830
rect 216 636 1026 671
rect 216 477 1026 512
rect 216 318 1026 353
rect 2700 216 2735 1026
rect 216 159 1026 194
rect 216 0 1026 35
rect 2859 216 2894 1026
rect 3018 216 3053 1026
rect 3177 216 3212 1026
rect 3336 216 3371 1026
rect 3495 216 3530 1026
rect 3654 216 3689 1026
rect 3813 216 3848 1026
rect 3972 216 4007 1026
rect 4131 216 4166 1026
<< locali >>
rect -75 1431 0 1466
rect 1125 1307 1142 1431
rect 100 1148 117 1272
rect 1125 989 1142 1113
rect 2735 1125 2859 1142
rect 3053 1125 3177 1142
rect 3371 1125 3495 1142
rect 3689 1125 3813 1142
rect 4007 1125 4131 1142
rect 100 830 117 954
rect 1125 671 1142 795
rect 100 512 117 636
rect 1125 353 1142 477
rect 100 194 117 318
rect 1125 35 1142 159
rect -75 0 0 35
rect 2894 100 3018 117
rect 3212 100 3336 117
rect 3530 100 3654 117
rect 3848 100 3972 117
rect 2700 -75 2735 0
rect 4131 -75 4166 0
<< end >>
