magic
tech sky130A
timestamp 1615384503
<< nwell >>
rect 954 1582 1097 9618
<< pmos >>
rect 1000 1600 1050 9600
<< pdiff >>
rect 972 1600 1000 9600
rect 1050 1600 1079 9600
<< poly >>
rect 1000 9600 1050 9625
rect 1000 1575 1050 1600
<< metal1 >>
rect 0 9700 29104 10000
rect 0 0 29104 500
<< properties >>
string FIXED_BBOX 0 0 29104 10000
<< end >>
